
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity project_tb is
end project_tb;

architecture projecttb of project_tb is
constant c_CLOCK_PERIOD         : time := 15 ns;
signal   tb_done                : std_logic;
signal   mem_address            : std_logic_vector (15 downto 0) := (others => '0');
signal   tb_rst                 : std_logic := '0';
signal   tb_start               : std_logic := '0';
signal   tb_clk                 : std_logic := '0';
signal   mem_o_data,mem_i_data  : std_logic_vector (7 downto 0);
signal   enable_wire            : std_logic;
signal   mem_we                 : std_logic;

type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);

signal i: std_logic_vector(1 downto 0) := "00";


signal RAM: ram_type := (0 => std_logic_vector(to_unsigned(42, 8)),
			1 => std_logic_vector(to_unsigned(41, 8)),
			2 => std_logic_vector(to_unsigned(141, 8)),
			3 => std_logic_vector(to_unsigned(168, 8)),
			4 => std_logic_vector(to_unsigned(3, 8)),
			5 => std_logic_vector(to_unsigned(72, 8)),
			6 => std_logic_vector(to_unsigned(22, 8)),
			7 => std_logic_vector(to_unsigned(220, 8)),
			8 => std_logic_vector(to_unsigned(224, 8)),
			9 => std_logic_vector(to_unsigned(54, 8)),
			10 => std_logic_vector(to_unsigned(97, 8)),
			11 => std_logic_vector(to_unsigned(12, 8)),
			12 => std_logic_vector(to_unsigned(148, 8)),
			13 => std_logic_vector(to_unsigned(10, 8)),
			14 => std_logic_vector(to_unsigned(41, 8)),
			15 => std_logic_vector(to_unsigned(50, 8)),
			16 => std_logic_vector(to_unsigned(142, 8)),
			17 => std_logic_vector(to_unsigned(252, 8)),
			18 => std_logic_vector(to_unsigned(143, 8)),
			19 => std_logic_vector(to_unsigned(203, 8)),
			20 => std_logic_vector(to_unsigned(33, 8)),
			21 => std_logic_vector(to_unsigned(82, 8)),
			22 => std_logic_vector(to_unsigned(112, 8)),
			23 => std_logic_vector(to_unsigned(241, 8)),
			24 => std_logic_vector(to_unsigned(159, 8)),
			25 => std_logic_vector(to_unsigned(47, 8)),
			26 => std_logic_vector(to_unsigned(50, 8)),
			27 => std_logic_vector(to_unsigned(73, 8)),
			28 => std_logic_vector(to_unsigned(140, 8)),
			29 => std_logic_vector(to_unsigned(121, 8)),
			30 => std_logic_vector(to_unsigned(204, 8)),
			31 => std_logic_vector(to_unsigned(216, 8)),
			32 => std_logic_vector(to_unsigned(200, 8)),
			33 => std_logic_vector(to_unsigned(181, 8)),
			34 => std_logic_vector(to_unsigned(109, 8)),
			35 => std_logic_vector(to_unsigned(174, 8)),
			36 => std_logic_vector(to_unsigned(200, 8)),
			37 => std_logic_vector(to_unsigned(105, 8)),
			38 => std_logic_vector(to_unsigned(157, 8)),
			39 => std_logic_vector(to_unsigned(108, 8)),
			40 => std_logic_vector(to_unsigned(207, 8)),
			41 => std_logic_vector(to_unsigned(64, 8)),
			42 => std_logic_vector(to_unsigned(60, 8)),
			43 => std_logic_vector(to_unsigned(242, 8)),
			44 => std_logic_vector(to_unsigned(17, 8)),
			45 => std_logic_vector(to_unsigned(170, 8)),
			46 => std_logic_vector(to_unsigned(245, 8)),
			47 => std_logic_vector(to_unsigned(106, 8)),
			48 => std_logic_vector(to_unsigned(201, 8)),
			49 => std_logic_vector(to_unsigned(120, 8)),
			50 => std_logic_vector(to_unsigned(90, 8)),
			51 => std_logic_vector(to_unsigned(107, 8)),
			52 => std_logic_vector(to_unsigned(249, 8)),
			53 => std_logic_vector(to_unsigned(12, 8)),
			54 => std_logic_vector(to_unsigned(176, 8)),
			55 => std_logic_vector(to_unsigned(170, 8)),
			56 => std_logic_vector(to_unsigned(249, 8)),
			57 => std_logic_vector(to_unsigned(188, 8)),
			58 => std_logic_vector(to_unsigned(86, 8)),
			59 => std_logic_vector(to_unsigned(37, 8)),
			60 => std_logic_vector(to_unsigned(83, 8)),
			61 => std_logic_vector(to_unsigned(172, 8)),
			62 => std_logic_vector(to_unsigned(208, 8)),
			63 => std_logic_vector(to_unsigned(214, 8)),
			64 => std_logic_vector(to_unsigned(35, 8)),
			65 => std_logic_vector(to_unsigned(122, 8)),
			66 => std_logic_vector(to_unsigned(217, 8)),
			67 => std_logic_vector(to_unsigned(154, 8)),
			68 => std_logic_vector(to_unsigned(187, 8)),
			69 => std_logic_vector(to_unsigned(130, 8)),
			70 => std_logic_vector(to_unsigned(115, 8)),
			71 => std_logic_vector(to_unsigned(218, 8)),
			72 => std_logic_vector(to_unsigned(180, 8)),
			73 => std_logic_vector(to_unsigned(127, 8)),
			74 => std_logic_vector(to_unsigned(48, 8)),
			75 => std_logic_vector(to_unsigned(112, 8)),
			76 => std_logic_vector(to_unsigned(47, 8)),
			77 => std_logic_vector(to_unsigned(213, 8)),
			78 => std_logic_vector(to_unsigned(127, 8)),
			79 => std_logic_vector(to_unsigned(120, 8)),
			80 => std_logic_vector(to_unsigned(193, 8)),
			81 => std_logic_vector(to_unsigned(143, 8)),
			82 => std_logic_vector(to_unsigned(151, 8)),
			83 => std_logic_vector(to_unsigned(5, 8)),
			84 => std_logic_vector(to_unsigned(111, 8)),
			85 => std_logic_vector(to_unsigned(29, 8)),
			86 => std_logic_vector(to_unsigned(124, 8)),
			87 => std_logic_vector(to_unsigned(35, 8)),
			88 => std_logic_vector(to_unsigned(192, 8)),
			89 => std_logic_vector(to_unsigned(129, 8)),
			90 => std_logic_vector(to_unsigned(227, 8)),
			91 => std_logic_vector(to_unsigned(108, 8)),
			92 => std_logic_vector(to_unsigned(164, 8)),
			93 => std_logic_vector(to_unsigned(0, 8)),
			94 => std_logic_vector(to_unsigned(158, 8)),
			95 => std_logic_vector(to_unsigned(188, 8)),
			96 => std_logic_vector(to_unsigned(108, 8)),
			97 => std_logic_vector(to_unsigned(81, 8)),
			98 => std_logic_vector(to_unsigned(98, 8)),
			99 => std_logic_vector(to_unsigned(144, 8)),
			100 => std_logic_vector(to_unsigned(14, 8)),
			101 => std_logic_vector(to_unsigned(203, 8)),
			102 => std_logic_vector(to_unsigned(205, 8)),
			103 => std_logic_vector(to_unsigned(59, 8)),
			104 => std_logic_vector(to_unsigned(220, 8)),
			105 => std_logic_vector(to_unsigned(217, 8)),
			106 => std_logic_vector(to_unsigned(147, 8)),
			107 => std_logic_vector(to_unsigned(128, 8)),
			108 => std_logic_vector(to_unsigned(219, 8)),
			109 => std_logic_vector(to_unsigned(65, 8)),
			110 => std_logic_vector(to_unsigned(95, 8)),
			111 => std_logic_vector(to_unsigned(64, 8)),
			112 => std_logic_vector(to_unsigned(228, 8)),
			113 => std_logic_vector(to_unsigned(144, 8)),
			114 => std_logic_vector(to_unsigned(118, 8)),
			115 => std_logic_vector(to_unsigned(157, 8)),
			116 => std_logic_vector(to_unsigned(97, 8)),
			117 => std_logic_vector(to_unsigned(246, 8)),
			118 => std_logic_vector(to_unsigned(36, 8)),
			119 => std_logic_vector(to_unsigned(43, 8)),
			120 => std_logic_vector(to_unsigned(251, 8)),
			121 => std_logic_vector(to_unsigned(120, 8)),
			122 => std_logic_vector(to_unsigned(125, 8)),
			123 => std_logic_vector(to_unsigned(100, 8)),
			124 => std_logic_vector(to_unsigned(97, 8)),
			125 => std_logic_vector(to_unsigned(71, 8)),
			126 => std_logic_vector(to_unsigned(7, 8)),
			127 => std_logic_vector(to_unsigned(17, 8)),
			128 => std_logic_vector(to_unsigned(112, 8)),
			129 => std_logic_vector(to_unsigned(93, 8)),
			130 => std_logic_vector(to_unsigned(196, 8)),
			131 => std_logic_vector(to_unsigned(191, 8)),
			132 => std_logic_vector(to_unsigned(146, 8)),
			133 => std_logic_vector(to_unsigned(104, 8)),
			134 => std_logic_vector(to_unsigned(61, 8)),
			135 => std_logic_vector(to_unsigned(49, 8)),
			136 => std_logic_vector(to_unsigned(136, 8)),
			137 => std_logic_vector(to_unsigned(233, 8)),
			138 => std_logic_vector(to_unsigned(100, 8)),
			139 => std_logic_vector(to_unsigned(40, 8)),
			140 => std_logic_vector(to_unsigned(153, 8)),
			141 => std_logic_vector(to_unsigned(92, 8)),
			142 => std_logic_vector(to_unsigned(207, 8)),
			143 => std_logic_vector(to_unsigned(27, 8)),
			144 => std_logic_vector(to_unsigned(156, 8)),
			145 => std_logic_vector(to_unsigned(105, 8)),
			146 => std_logic_vector(to_unsigned(75, 8)),
			147 => std_logic_vector(to_unsigned(80, 8)),
			148 => std_logic_vector(to_unsigned(220, 8)),
			149 => std_logic_vector(to_unsigned(3, 8)),
			150 => std_logic_vector(to_unsigned(90, 8)),
			151 => std_logic_vector(to_unsigned(119, 8)),
			152 => std_logic_vector(to_unsigned(195, 8)),
			153 => std_logic_vector(to_unsigned(62, 8)),
			154 => std_logic_vector(to_unsigned(83, 8)),
			155 => std_logic_vector(to_unsigned(124, 8)),
			156 => std_logic_vector(to_unsigned(14, 8)),
			157 => std_logic_vector(to_unsigned(102, 8)),
			158 => std_logic_vector(to_unsigned(247, 8)),
			159 => std_logic_vector(to_unsigned(217, 8)),
			160 => std_logic_vector(to_unsigned(126, 8)),
			161 => std_logic_vector(to_unsigned(201, 8)),
			162 => std_logic_vector(to_unsigned(193, 8)),
			163 => std_logic_vector(to_unsigned(142, 8)),
			164 => std_logic_vector(to_unsigned(183, 8)),
			165 => std_logic_vector(to_unsigned(4, 8)),
			166 => std_logic_vector(to_unsigned(69, 8)),
			167 => std_logic_vector(to_unsigned(98, 8)),
			168 => std_logic_vector(to_unsigned(85, 8)),
			169 => std_logic_vector(to_unsigned(51, 8)),
			170 => std_logic_vector(to_unsigned(88, 8)),
			171 => std_logic_vector(to_unsigned(50, 8)),
			172 => std_logic_vector(to_unsigned(72, 8)),
			173 => std_logic_vector(to_unsigned(235, 8)),
			174 => std_logic_vector(to_unsigned(211, 8)),
			175 => std_logic_vector(to_unsigned(5, 8)),
			176 => std_logic_vector(to_unsigned(203, 8)),
			177 => std_logic_vector(to_unsigned(217, 8)),
			178 => std_logic_vector(to_unsigned(172, 8)),
			179 => std_logic_vector(to_unsigned(214, 8)),
			180 => std_logic_vector(to_unsigned(134, 8)),
			181 => std_logic_vector(to_unsigned(113, 8)),
			182 => std_logic_vector(to_unsigned(80, 8)),
			183 => std_logic_vector(to_unsigned(16, 8)),
			184 => std_logic_vector(to_unsigned(211, 8)),
			185 => std_logic_vector(to_unsigned(26, 8)),
			186 => std_logic_vector(to_unsigned(97, 8)),
			187 => std_logic_vector(to_unsigned(87, 8)),
			188 => std_logic_vector(to_unsigned(204, 8)),
			189 => std_logic_vector(to_unsigned(113, 8)),
			190 => std_logic_vector(to_unsigned(28, 8)),
			191 => std_logic_vector(to_unsigned(185, 8)),
			192 => std_logic_vector(to_unsigned(200, 8)),
			193 => std_logic_vector(to_unsigned(92, 8)),
			194 => std_logic_vector(to_unsigned(87, 8)),
			195 => std_logic_vector(to_unsigned(38, 8)),
			196 => std_logic_vector(to_unsigned(121, 8)),
			197 => std_logic_vector(to_unsigned(181, 8)),
			198 => std_logic_vector(to_unsigned(4, 8)),
			199 => std_logic_vector(to_unsigned(1, 8)),
			200 => std_logic_vector(to_unsigned(130, 8)),
			201 => std_logic_vector(to_unsigned(172, 8)),
			202 => std_logic_vector(to_unsigned(136, 8)),
			203 => std_logic_vector(to_unsigned(196, 8)),
			204 => std_logic_vector(to_unsigned(134, 8)),
			205 => std_logic_vector(to_unsigned(66, 8)),
			206 => std_logic_vector(to_unsigned(102, 8)),
			207 => std_logic_vector(to_unsigned(52, 8)),
			208 => std_logic_vector(to_unsigned(143, 8)),
			209 => std_logic_vector(to_unsigned(88, 8)),
			210 => std_logic_vector(to_unsigned(184, 8)),
			211 => std_logic_vector(to_unsigned(212, 8)),
			212 => std_logic_vector(to_unsigned(245, 8)),
			213 => std_logic_vector(to_unsigned(120, 8)),
			214 => std_logic_vector(to_unsigned(5, 8)),
			215 => std_logic_vector(to_unsigned(247, 8)),
			216 => std_logic_vector(to_unsigned(62, 8)),
			217 => std_logic_vector(to_unsigned(209, 8)),
			218 => std_logic_vector(to_unsigned(204, 8)),
			219 => std_logic_vector(to_unsigned(139, 8)),
			220 => std_logic_vector(to_unsigned(191, 8)),
			221 => std_logic_vector(to_unsigned(135, 8)),
			222 => std_logic_vector(to_unsigned(229, 8)),
			223 => std_logic_vector(to_unsigned(105, 8)),
			224 => std_logic_vector(to_unsigned(162, 8)),
			225 => std_logic_vector(to_unsigned(141, 8)),
			226 => std_logic_vector(to_unsigned(20, 8)),
			227 => std_logic_vector(to_unsigned(160, 8)),
			228 => std_logic_vector(to_unsigned(25, 8)),
			229 => std_logic_vector(to_unsigned(143, 8)),
			230 => std_logic_vector(to_unsigned(172, 8)),
			231 => std_logic_vector(to_unsigned(77, 8)),
			232 => std_logic_vector(to_unsigned(239, 8)),
			233 => std_logic_vector(to_unsigned(185, 8)),
			234 => std_logic_vector(to_unsigned(183, 8)),
			235 => std_logic_vector(to_unsigned(185, 8)),
			236 => std_logic_vector(to_unsigned(120, 8)),
			237 => std_logic_vector(to_unsigned(62, 8)),
			238 => std_logic_vector(to_unsigned(157, 8)),
			239 => std_logic_vector(to_unsigned(126, 8)),
			240 => std_logic_vector(to_unsigned(147, 8)),
			241 => std_logic_vector(to_unsigned(43, 8)),
			242 => std_logic_vector(to_unsigned(169, 8)),
			243 => std_logic_vector(to_unsigned(82, 8)),
			244 => std_logic_vector(to_unsigned(122, 8)),
			245 => std_logic_vector(to_unsigned(119, 8)),
			246 => std_logic_vector(to_unsigned(117, 8)),
			247 => std_logic_vector(to_unsigned(25, 8)),
			248 => std_logic_vector(to_unsigned(25, 8)),
			249 => std_logic_vector(to_unsigned(129, 8)),
			250 => std_logic_vector(to_unsigned(219, 8)),
			251 => std_logic_vector(to_unsigned(163, 8)),
			252 => std_logic_vector(to_unsigned(57, 8)),
			253 => std_logic_vector(to_unsigned(238, 8)),
			254 => std_logic_vector(to_unsigned(210, 8)),
			255 => std_logic_vector(to_unsigned(129, 8)),
			256 => std_logic_vector(to_unsigned(148, 8)),
			257 => std_logic_vector(to_unsigned(74, 8)),
			258 => std_logic_vector(to_unsigned(165, 8)),
			259 => std_logic_vector(to_unsigned(121, 8)),
			260 => std_logic_vector(to_unsigned(7, 8)),
			261 => std_logic_vector(to_unsigned(35, 8)),
			262 => std_logic_vector(to_unsigned(22, 8)),
			263 => std_logic_vector(to_unsigned(136, 8)),
			264 => std_logic_vector(to_unsigned(209, 8)),
			265 => std_logic_vector(to_unsigned(65, 8)),
			266 => std_logic_vector(to_unsigned(119, 8)),
			267 => std_logic_vector(to_unsigned(222, 8)),
			268 => std_logic_vector(to_unsigned(237, 8)),
			269 => std_logic_vector(to_unsigned(90, 8)),
			270 => std_logic_vector(to_unsigned(26, 8)),
			271 => std_logic_vector(to_unsigned(246, 8)),
			272 => std_logic_vector(to_unsigned(103, 8)),
			273 => std_logic_vector(to_unsigned(229, 8)),
			274 => std_logic_vector(to_unsigned(187, 8)),
			275 => std_logic_vector(to_unsigned(192, 8)),
			276 => std_logic_vector(to_unsigned(36, 8)),
			277 => std_logic_vector(to_unsigned(109, 8)),
			278 => std_logic_vector(to_unsigned(164, 8)),
			279 => std_logic_vector(to_unsigned(173, 8)),
			280 => std_logic_vector(to_unsigned(54, 8)),
			281 => std_logic_vector(to_unsigned(250, 8)),
			282 => std_logic_vector(to_unsigned(184, 8)),
			283 => std_logic_vector(to_unsigned(145, 8)),
			284 => std_logic_vector(to_unsigned(180, 8)),
			285 => std_logic_vector(to_unsigned(46, 8)),
			286 => std_logic_vector(to_unsigned(237, 8)),
			287 => std_logic_vector(to_unsigned(233, 8)),
			288 => std_logic_vector(to_unsigned(49, 8)),
			289 => std_logic_vector(to_unsigned(110, 8)),
			290 => std_logic_vector(to_unsigned(133, 8)),
			291 => std_logic_vector(to_unsigned(247, 8)),
			292 => std_logic_vector(to_unsigned(121, 8)),
			293 => std_logic_vector(to_unsigned(39, 8)),
			294 => std_logic_vector(to_unsigned(58, 8)),
			295 => std_logic_vector(to_unsigned(250, 8)),
			296 => std_logic_vector(to_unsigned(151, 8)),
			297 => std_logic_vector(to_unsigned(6, 8)),
			298 => std_logic_vector(to_unsigned(232, 8)),
			299 => std_logic_vector(to_unsigned(170, 8)),
			300 => std_logic_vector(to_unsigned(255, 8)),
			301 => std_logic_vector(to_unsigned(116, 8)),
			302 => std_logic_vector(to_unsigned(169, 8)),
			303 => std_logic_vector(to_unsigned(60, 8)),
			304 => std_logic_vector(to_unsigned(8, 8)),
			305 => std_logic_vector(to_unsigned(245, 8)),
			306 => std_logic_vector(to_unsigned(91, 8)),
			307 => std_logic_vector(to_unsigned(236, 8)),
			308 => std_logic_vector(to_unsigned(14, 8)),
			309 => std_logic_vector(to_unsigned(83, 8)),
			310 => std_logic_vector(to_unsigned(70, 8)),
			311 => std_logic_vector(to_unsigned(224, 8)),
			312 => std_logic_vector(to_unsigned(139, 8)),
			313 => std_logic_vector(to_unsigned(116, 8)),
			314 => std_logic_vector(to_unsigned(163, 8)),
			315 => std_logic_vector(to_unsigned(33, 8)),
			316 => std_logic_vector(to_unsigned(38, 8)),
			317 => std_logic_vector(to_unsigned(114, 8)),
			318 => std_logic_vector(to_unsigned(111, 8)),
			319 => std_logic_vector(to_unsigned(94, 8)),
			320 => std_logic_vector(to_unsigned(89, 8)),
			321 => std_logic_vector(to_unsigned(143, 8)),
			322 => std_logic_vector(to_unsigned(59, 8)),
			323 => std_logic_vector(to_unsigned(229, 8)),
			324 => std_logic_vector(to_unsigned(245, 8)),
			325 => std_logic_vector(to_unsigned(99, 8)),
			326 => std_logic_vector(to_unsigned(85, 8)),
			327 => std_logic_vector(to_unsigned(234, 8)),
			328 => std_logic_vector(to_unsigned(17, 8)),
			329 => std_logic_vector(to_unsigned(0, 8)),
			330 => std_logic_vector(to_unsigned(198, 8)),
			331 => std_logic_vector(to_unsigned(176, 8)),
			332 => std_logic_vector(to_unsigned(192, 8)),
			333 => std_logic_vector(to_unsigned(226, 8)),
			334 => std_logic_vector(to_unsigned(78, 8)),
			335 => std_logic_vector(to_unsigned(113, 8)),
			336 => std_logic_vector(to_unsigned(85, 8)),
			337 => std_logic_vector(to_unsigned(74, 8)),
			338 => std_logic_vector(to_unsigned(202, 8)),
			339 => std_logic_vector(to_unsigned(106, 8)),
			340 => std_logic_vector(to_unsigned(91, 8)),
			341 => std_logic_vector(to_unsigned(41, 8)),
			342 => std_logic_vector(to_unsigned(107, 8)),
			343 => std_logic_vector(to_unsigned(27, 8)),
			344 => std_logic_vector(to_unsigned(120, 8)),
			345 => std_logic_vector(to_unsigned(227, 8)),
			346 => std_logic_vector(to_unsigned(41, 8)),
			347 => std_logic_vector(to_unsigned(50, 8)),
			348 => std_logic_vector(to_unsigned(15, 8)),
			349 => std_logic_vector(to_unsigned(124, 8)),
			350 => std_logic_vector(to_unsigned(129, 8)),
			351 => std_logic_vector(to_unsigned(123, 8)),
			352 => std_logic_vector(to_unsigned(21, 8)),
			353 => std_logic_vector(to_unsigned(227, 8)),
			354 => std_logic_vector(to_unsigned(61, 8)),
			355 => std_logic_vector(to_unsigned(51, 8)),
			356 => std_logic_vector(to_unsigned(61, 8)),
			357 => std_logic_vector(to_unsigned(245, 8)),
			358 => std_logic_vector(to_unsigned(0, 8)),
			359 => std_logic_vector(to_unsigned(142, 8)),
			360 => std_logic_vector(to_unsigned(172, 8)),
			361 => std_logic_vector(to_unsigned(232, 8)),
			362 => std_logic_vector(to_unsigned(213, 8)),
			363 => std_logic_vector(to_unsigned(199, 8)),
			364 => std_logic_vector(to_unsigned(12, 8)),
			365 => std_logic_vector(to_unsigned(174, 8)),
			366 => std_logic_vector(to_unsigned(26, 8)),
			367 => std_logic_vector(to_unsigned(131, 8)),
			368 => std_logic_vector(to_unsigned(245, 8)),
			369 => std_logic_vector(to_unsigned(104, 8)),
			370 => std_logic_vector(to_unsigned(48, 8)),
			371 => std_logic_vector(to_unsigned(62, 8)),
			372 => std_logic_vector(to_unsigned(252, 8)),
			373 => std_logic_vector(to_unsigned(188, 8)),
			374 => std_logic_vector(to_unsigned(233, 8)),
			375 => std_logic_vector(to_unsigned(87, 8)),
			376 => std_logic_vector(to_unsigned(240, 8)),
			377 => std_logic_vector(to_unsigned(209, 8)),
			378 => std_logic_vector(to_unsigned(156, 8)),
			379 => std_logic_vector(to_unsigned(94, 8)),
			380 => std_logic_vector(to_unsigned(112, 8)),
			381 => std_logic_vector(to_unsigned(176, 8)),
			382 => std_logic_vector(to_unsigned(202, 8)),
			383 => std_logic_vector(to_unsigned(10, 8)),
			384 => std_logic_vector(to_unsigned(172, 8)),
			385 => std_logic_vector(to_unsigned(0, 8)),
			386 => std_logic_vector(to_unsigned(147, 8)),
			387 => std_logic_vector(to_unsigned(99, 8)),
			388 => std_logic_vector(to_unsigned(23, 8)),
			389 => std_logic_vector(to_unsigned(126, 8)),
			390 => std_logic_vector(to_unsigned(96, 8)),
			391 => std_logic_vector(to_unsigned(24, 8)),
			392 => std_logic_vector(to_unsigned(8, 8)),
			393 => std_logic_vector(to_unsigned(106, 8)),
			394 => std_logic_vector(to_unsigned(112, 8)),
			395 => std_logic_vector(to_unsigned(200, 8)),
			396 => std_logic_vector(to_unsigned(28, 8)),
			397 => std_logic_vector(to_unsigned(214, 8)),
			398 => std_logic_vector(to_unsigned(178, 8)),
			399 => std_logic_vector(to_unsigned(184, 8)),
			400 => std_logic_vector(to_unsigned(204, 8)),
			401 => std_logic_vector(to_unsigned(149, 8)),
			402 => std_logic_vector(to_unsigned(238, 8)),
			403 => std_logic_vector(to_unsigned(229, 8)),
			404 => std_logic_vector(to_unsigned(102, 8)),
			405 => std_logic_vector(to_unsigned(21, 8)),
			406 => std_logic_vector(to_unsigned(201, 8)),
			407 => std_logic_vector(to_unsigned(161, 8)),
			408 => std_logic_vector(to_unsigned(32, 8)),
			409 => std_logic_vector(to_unsigned(219, 8)),
			410 => std_logic_vector(to_unsigned(154, 8)),
			411 => std_logic_vector(to_unsigned(29, 8)),
			412 => std_logic_vector(to_unsigned(22, 8)),
			413 => std_logic_vector(to_unsigned(86, 8)),
			414 => std_logic_vector(to_unsigned(160, 8)),
			415 => std_logic_vector(to_unsigned(147, 8)),
			416 => std_logic_vector(to_unsigned(220, 8)),
			417 => std_logic_vector(to_unsigned(152, 8)),
			418 => std_logic_vector(to_unsigned(174, 8)),
			419 => std_logic_vector(to_unsigned(162, 8)),
			420 => std_logic_vector(to_unsigned(100, 8)),
			421 => std_logic_vector(to_unsigned(174, 8)),
			422 => std_logic_vector(to_unsigned(9, 8)),
			423 => std_logic_vector(to_unsigned(160, 8)),
			424 => std_logic_vector(to_unsigned(177, 8)),
			425 => std_logic_vector(to_unsigned(36, 8)),
			426 => std_logic_vector(to_unsigned(184, 8)),
			427 => std_logic_vector(to_unsigned(128, 8)),
			428 => std_logic_vector(to_unsigned(216, 8)),
			429 => std_logic_vector(to_unsigned(33, 8)),
			430 => std_logic_vector(to_unsigned(68, 8)),
			431 => std_logic_vector(to_unsigned(183, 8)),
			432 => std_logic_vector(to_unsigned(122, 8)),
			433 => std_logic_vector(to_unsigned(20, 8)),
			434 => std_logic_vector(to_unsigned(64, 8)),
			435 => std_logic_vector(to_unsigned(161, 8)),
			436 => std_logic_vector(to_unsigned(8, 8)),
			437 => std_logic_vector(to_unsigned(165, 8)),
			438 => std_logic_vector(to_unsigned(139, 8)),
			439 => std_logic_vector(to_unsigned(212, 8)),
			440 => std_logic_vector(to_unsigned(225, 8)),
			441 => std_logic_vector(to_unsigned(26, 8)),
			442 => std_logic_vector(to_unsigned(245, 8)),
			443 => std_logic_vector(to_unsigned(240, 8)),
			444 => std_logic_vector(to_unsigned(6, 8)),
			445 => std_logic_vector(to_unsigned(127, 8)),
			446 => std_logic_vector(to_unsigned(80, 8)),
			447 => std_logic_vector(to_unsigned(185, 8)),
			448 => std_logic_vector(to_unsigned(15, 8)),
			449 => std_logic_vector(to_unsigned(33, 8)),
			450 => std_logic_vector(to_unsigned(50, 8)),
			451 => std_logic_vector(to_unsigned(108, 8)),
			452 => std_logic_vector(to_unsigned(131, 8)),
			453 => std_logic_vector(to_unsigned(16, 8)),
			454 => std_logic_vector(to_unsigned(36, 8)),
			455 => std_logic_vector(to_unsigned(209, 8)),
			456 => std_logic_vector(to_unsigned(87, 8)),
			457 => std_logic_vector(to_unsigned(83, 8)),
			458 => std_logic_vector(to_unsigned(111, 8)),
			459 => std_logic_vector(to_unsigned(227, 8)),
			460 => std_logic_vector(to_unsigned(47, 8)),
			461 => std_logic_vector(to_unsigned(124, 8)),
			462 => std_logic_vector(to_unsigned(124, 8)),
			463 => std_logic_vector(to_unsigned(152, 8)),
			464 => std_logic_vector(to_unsigned(98, 8)),
			465 => std_logic_vector(to_unsigned(109, 8)),
			466 => std_logic_vector(to_unsigned(98, 8)),
			467 => std_logic_vector(to_unsigned(11, 8)),
			468 => std_logic_vector(to_unsigned(161, 8)),
			469 => std_logic_vector(to_unsigned(125, 8)),
			470 => std_logic_vector(to_unsigned(31, 8)),
			471 => std_logic_vector(to_unsigned(199, 8)),
			472 => std_logic_vector(to_unsigned(124, 8)),
			473 => std_logic_vector(to_unsigned(85, 8)),
			474 => std_logic_vector(to_unsigned(24, 8)),
			475 => std_logic_vector(to_unsigned(246, 8)),
			476 => std_logic_vector(to_unsigned(142, 8)),
			477 => std_logic_vector(to_unsigned(39, 8)),
			478 => std_logic_vector(to_unsigned(166, 8)),
			479 => std_logic_vector(to_unsigned(136, 8)),
			480 => std_logic_vector(to_unsigned(180, 8)),
			481 => std_logic_vector(to_unsigned(71, 8)),
			482 => std_logic_vector(to_unsigned(64, 8)),
			483 => std_logic_vector(to_unsigned(90, 8)),
			484 => std_logic_vector(to_unsigned(61, 8)),
			485 => std_logic_vector(to_unsigned(245, 8)),
			486 => std_logic_vector(to_unsigned(251, 8)),
			487 => std_logic_vector(to_unsigned(203, 8)),
			488 => std_logic_vector(to_unsigned(62, 8)),
			489 => std_logic_vector(to_unsigned(24, 8)),
			490 => std_logic_vector(to_unsigned(31, 8)),
			491 => std_logic_vector(to_unsigned(101, 8)),
			492 => std_logic_vector(to_unsigned(21, 8)),
			493 => std_logic_vector(to_unsigned(37, 8)),
			494 => std_logic_vector(to_unsigned(245, 8)),
			495 => std_logic_vector(to_unsigned(216, 8)),
			496 => std_logic_vector(to_unsigned(133, 8)),
			497 => std_logic_vector(to_unsigned(90, 8)),
			498 => std_logic_vector(to_unsigned(181, 8)),
			499 => std_logic_vector(to_unsigned(173, 8)),
			500 => std_logic_vector(to_unsigned(98, 8)),
			501 => std_logic_vector(to_unsigned(132, 8)),
			502 => std_logic_vector(to_unsigned(118, 8)),
			503 => std_logic_vector(to_unsigned(116, 8)),
			504 => std_logic_vector(to_unsigned(200, 8)),
			505 => std_logic_vector(to_unsigned(6, 8)),
			506 => std_logic_vector(to_unsigned(92, 8)),
			507 => std_logic_vector(to_unsigned(123, 8)),
			508 => std_logic_vector(to_unsigned(159, 8)),
			509 => std_logic_vector(to_unsigned(20, 8)),
			510 => std_logic_vector(to_unsigned(62, 8)),
			511 => std_logic_vector(to_unsigned(146, 8)),
			512 => std_logic_vector(to_unsigned(36, 8)),
			513 => std_logic_vector(to_unsigned(44, 8)),
			514 => std_logic_vector(to_unsigned(8, 8)),
			515 => std_logic_vector(to_unsigned(70, 8)),
			516 => std_logic_vector(to_unsigned(152, 8)),
			517 => std_logic_vector(to_unsigned(250, 8)),
			518 => std_logic_vector(to_unsigned(85, 8)),
			519 => std_logic_vector(to_unsigned(183, 8)),
			520 => std_logic_vector(to_unsigned(141, 8)),
			521 => std_logic_vector(to_unsigned(206, 8)),
			522 => std_logic_vector(to_unsigned(81, 8)),
			523 => std_logic_vector(to_unsigned(187, 8)),
			524 => std_logic_vector(to_unsigned(249, 8)),
			525 => std_logic_vector(to_unsigned(203, 8)),
			526 => std_logic_vector(to_unsigned(91, 8)),
			527 => std_logic_vector(to_unsigned(55, 8)),
			528 => std_logic_vector(to_unsigned(70, 8)),
			529 => std_logic_vector(to_unsigned(65, 8)),
			530 => std_logic_vector(to_unsigned(150, 8)),
			531 => std_logic_vector(to_unsigned(131, 8)),
			532 => std_logic_vector(to_unsigned(101, 8)),
			533 => std_logic_vector(to_unsigned(11, 8)),
			534 => std_logic_vector(to_unsigned(19, 8)),
			535 => std_logic_vector(to_unsigned(74, 8)),
			536 => std_logic_vector(to_unsigned(180, 8)),
			537 => std_logic_vector(to_unsigned(1, 8)),
			538 => std_logic_vector(to_unsigned(18, 8)),
			539 => std_logic_vector(to_unsigned(128, 8)),
			540 => std_logic_vector(to_unsigned(127, 8)),
			541 => std_logic_vector(to_unsigned(156, 8)),
			542 => std_logic_vector(to_unsigned(109, 8)),
			543 => std_logic_vector(to_unsigned(242, 8)),
			544 => std_logic_vector(to_unsigned(207, 8)),
			545 => std_logic_vector(to_unsigned(164, 8)),
			546 => std_logic_vector(to_unsigned(173, 8)),
			547 => std_logic_vector(to_unsigned(72, 8)),
			548 => std_logic_vector(to_unsigned(128, 8)),
			549 => std_logic_vector(to_unsigned(122, 8)),
			550 => std_logic_vector(to_unsigned(214, 8)),
			551 => std_logic_vector(to_unsigned(182, 8)),
			552 => std_logic_vector(to_unsigned(6, 8)),
			553 => std_logic_vector(to_unsigned(173, 8)),
			554 => std_logic_vector(to_unsigned(80, 8)),
			555 => std_logic_vector(to_unsigned(1, 8)),
			556 => std_logic_vector(to_unsigned(188, 8)),
			557 => std_logic_vector(to_unsigned(187, 8)),
			558 => std_logic_vector(to_unsigned(124, 8)),
			559 => std_logic_vector(to_unsigned(74, 8)),
			560 => std_logic_vector(to_unsigned(21, 8)),
			561 => std_logic_vector(to_unsigned(189, 8)),
			562 => std_logic_vector(to_unsigned(178, 8)),
			563 => std_logic_vector(to_unsigned(231, 8)),
			564 => std_logic_vector(to_unsigned(12, 8)),
			565 => std_logic_vector(to_unsigned(17, 8)),
			566 => std_logic_vector(to_unsigned(112, 8)),
			567 => std_logic_vector(to_unsigned(56, 8)),
			568 => std_logic_vector(to_unsigned(229, 8)),
			569 => std_logic_vector(to_unsigned(205, 8)),
			570 => std_logic_vector(to_unsigned(61, 8)),
			571 => std_logic_vector(to_unsigned(201, 8)),
			572 => std_logic_vector(to_unsigned(137, 8)),
			573 => std_logic_vector(to_unsigned(100, 8)),
			574 => std_logic_vector(to_unsigned(60, 8)),
			575 => std_logic_vector(to_unsigned(11, 8)),
			576 => std_logic_vector(to_unsigned(200, 8)),
			577 => std_logic_vector(to_unsigned(163, 8)),
			578 => std_logic_vector(to_unsigned(66, 8)),
			579 => std_logic_vector(to_unsigned(31, 8)),
			580 => std_logic_vector(to_unsigned(159, 8)),
			581 => std_logic_vector(to_unsigned(255, 8)),
			582 => std_logic_vector(to_unsigned(178, 8)),
			583 => std_logic_vector(to_unsigned(248, 8)),
			584 => std_logic_vector(to_unsigned(159, 8)),
			585 => std_logic_vector(to_unsigned(179, 8)),
			586 => std_logic_vector(to_unsigned(182, 8)),
			587 => std_logic_vector(to_unsigned(40, 8)),
			588 => std_logic_vector(to_unsigned(175, 8)),
			589 => std_logic_vector(to_unsigned(183, 8)),
			590 => std_logic_vector(to_unsigned(146, 8)),
			591 => std_logic_vector(to_unsigned(52, 8)),
			592 => std_logic_vector(to_unsigned(45, 8)),
			593 => std_logic_vector(to_unsigned(102, 8)),
			594 => std_logic_vector(to_unsigned(51, 8)),
			595 => std_logic_vector(to_unsigned(71, 8)),
			596 => std_logic_vector(to_unsigned(86, 8)),
			597 => std_logic_vector(to_unsigned(119, 8)),
			598 => std_logic_vector(to_unsigned(192, 8)),
			599 => std_logic_vector(to_unsigned(12, 8)),
			600 => std_logic_vector(to_unsigned(6, 8)),
			601 => std_logic_vector(to_unsigned(191, 8)),
			602 => std_logic_vector(to_unsigned(115, 8)),
			603 => std_logic_vector(to_unsigned(15, 8)),
			604 => std_logic_vector(to_unsigned(95, 8)),
			605 => std_logic_vector(to_unsigned(189, 8)),
			606 => std_logic_vector(to_unsigned(102, 8)),
			607 => std_logic_vector(to_unsigned(87, 8)),
			608 => std_logic_vector(to_unsigned(150, 8)),
			609 => std_logic_vector(to_unsigned(187, 8)),
			610 => std_logic_vector(to_unsigned(255, 8)),
			611 => std_logic_vector(to_unsigned(95, 8)),
			612 => std_logic_vector(to_unsigned(230, 8)),
			613 => std_logic_vector(to_unsigned(94, 8)),
			614 => std_logic_vector(to_unsigned(66, 8)),
			615 => std_logic_vector(to_unsigned(219, 8)),
			616 => std_logic_vector(to_unsigned(82, 8)),
			617 => std_logic_vector(to_unsigned(151, 8)),
			618 => std_logic_vector(to_unsigned(172, 8)),
			619 => std_logic_vector(to_unsigned(191, 8)),
			620 => std_logic_vector(to_unsigned(213, 8)),
			621 => std_logic_vector(to_unsigned(152, 8)),
			622 => std_logic_vector(to_unsigned(77, 8)),
			623 => std_logic_vector(to_unsigned(29, 8)),
			624 => std_logic_vector(to_unsigned(11, 8)),
			625 => std_logic_vector(to_unsigned(220, 8)),
			626 => std_logic_vector(to_unsigned(196, 8)),
			627 => std_logic_vector(to_unsigned(175, 8)),
			628 => std_logic_vector(to_unsigned(100, 8)),
			629 => std_logic_vector(to_unsigned(63, 8)),
			630 => std_logic_vector(to_unsigned(14, 8)),
			631 => std_logic_vector(to_unsigned(231, 8)),
			632 => std_logic_vector(to_unsigned(117, 8)),
			633 => std_logic_vector(to_unsigned(5, 8)),
			634 => std_logic_vector(to_unsigned(223, 8)),
			635 => std_logic_vector(to_unsigned(35, 8)),
			636 => std_logic_vector(to_unsigned(189, 8)),
			637 => std_logic_vector(to_unsigned(192, 8)),
			638 => std_logic_vector(to_unsigned(155, 8)),
			639 => std_logic_vector(to_unsigned(195, 8)),
			640 => std_logic_vector(to_unsigned(11, 8)),
			641 => std_logic_vector(to_unsigned(247, 8)),
			642 => std_logic_vector(to_unsigned(66, 8)),
			643 => std_logic_vector(to_unsigned(118, 8)),
			644 => std_logic_vector(to_unsigned(211, 8)),
			645 => std_logic_vector(to_unsigned(37, 8)),
			646 => std_logic_vector(to_unsigned(32, 8)),
			647 => std_logic_vector(to_unsigned(184, 8)),
			648 => std_logic_vector(to_unsigned(193, 8)),
			649 => std_logic_vector(to_unsigned(106, 8)),
			650 => std_logic_vector(to_unsigned(102, 8)),
			651 => std_logic_vector(to_unsigned(224, 8)),
			652 => std_logic_vector(to_unsigned(103, 8)),
			653 => std_logic_vector(to_unsigned(18, 8)),
			654 => std_logic_vector(to_unsigned(61, 8)),
			655 => std_logic_vector(to_unsigned(129, 8)),
			656 => std_logic_vector(to_unsigned(63, 8)),
			657 => std_logic_vector(to_unsigned(76, 8)),
			658 => std_logic_vector(to_unsigned(195, 8)),
			659 => std_logic_vector(to_unsigned(200, 8)),
			660 => std_logic_vector(to_unsigned(163, 8)),
			661 => std_logic_vector(to_unsigned(55, 8)),
			662 => std_logic_vector(to_unsigned(50, 8)),
			663 => std_logic_vector(to_unsigned(205, 8)),
			664 => std_logic_vector(to_unsigned(143, 8)),
			665 => std_logic_vector(to_unsigned(152, 8)),
			666 => std_logic_vector(to_unsigned(224, 8)),
			667 => std_logic_vector(to_unsigned(239, 8)),
			668 => std_logic_vector(to_unsigned(163, 8)),
			669 => std_logic_vector(to_unsigned(208, 8)),
			670 => std_logic_vector(to_unsigned(93, 8)),
			671 => std_logic_vector(to_unsigned(226, 8)),
			672 => std_logic_vector(to_unsigned(220, 8)),
			673 => std_logic_vector(to_unsigned(235, 8)),
			674 => std_logic_vector(to_unsigned(242, 8)),
			675 => std_logic_vector(to_unsigned(18, 8)),
			676 => std_logic_vector(to_unsigned(104, 8)),
			677 => std_logic_vector(to_unsigned(255, 8)),
			678 => std_logic_vector(to_unsigned(206, 8)),
			679 => std_logic_vector(to_unsigned(184, 8)),
			680 => std_logic_vector(to_unsigned(76, 8)),
			681 => std_logic_vector(to_unsigned(211, 8)),
			682 => std_logic_vector(to_unsigned(77, 8)),
			683 => std_logic_vector(to_unsigned(19, 8)),
			684 => std_logic_vector(to_unsigned(246, 8)),
			685 => std_logic_vector(to_unsigned(3, 8)),
			686 => std_logic_vector(to_unsigned(31, 8)),
			687 => std_logic_vector(to_unsigned(14, 8)),
			688 => std_logic_vector(to_unsigned(158, 8)),
			689 => std_logic_vector(to_unsigned(113, 8)),
			690 => std_logic_vector(to_unsigned(141, 8)),
			691 => std_logic_vector(to_unsigned(133, 8)),
			692 => std_logic_vector(to_unsigned(110, 8)),
			693 => std_logic_vector(to_unsigned(202, 8)),
			694 => std_logic_vector(to_unsigned(145, 8)),
			695 => std_logic_vector(to_unsigned(210, 8)),
			696 => std_logic_vector(to_unsigned(146, 8)),
			697 => std_logic_vector(to_unsigned(64, 8)),
			698 => std_logic_vector(to_unsigned(146, 8)),
			699 => std_logic_vector(to_unsigned(247, 8)),
			700 => std_logic_vector(to_unsigned(226, 8)),
			701 => std_logic_vector(to_unsigned(130, 8)),
			702 => std_logic_vector(to_unsigned(46, 8)),
			703 => std_logic_vector(to_unsigned(236, 8)),
			704 => std_logic_vector(to_unsigned(207, 8)),
			705 => std_logic_vector(to_unsigned(126, 8)),
			706 => std_logic_vector(to_unsigned(21, 8)),
			707 => std_logic_vector(to_unsigned(202, 8)),
			708 => std_logic_vector(to_unsigned(182, 8)),
			709 => std_logic_vector(to_unsigned(26, 8)),
			710 => std_logic_vector(to_unsigned(150, 8)),
			711 => std_logic_vector(to_unsigned(233, 8)),
			712 => std_logic_vector(to_unsigned(21, 8)),
			713 => std_logic_vector(to_unsigned(41, 8)),
			714 => std_logic_vector(to_unsigned(165, 8)),
			715 => std_logic_vector(to_unsigned(72, 8)),
			716 => std_logic_vector(to_unsigned(202, 8)),
			717 => std_logic_vector(to_unsigned(200, 8)),
			718 => std_logic_vector(to_unsigned(158, 8)),
			719 => std_logic_vector(to_unsigned(60, 8)),
			720 => std_logic_vector(to_unsigned(126, 8)),
			721 => std_logic_vector(to_unsigned(22, 8)),
			722 => std_logic_vector(to_unsigned(136, 8)),
			723 => std_logic_vector(to_unsigned(118, 8)),
			724 => std_logic_vector(to_unsigned(17, 8)),
			725 => std_logic_vector(to_unsigned(182, 8)),
			726 => std_logic_vector(to_unsigned(230, 8)),
			727 => std_logic_vector(to_unsigned(86, 8)),
			728 => std_logic_vector(to_unsigned(25, 8)),
			729 => std_logic_vector(to_unsigned(129, 8)),
			730 => std_logic_vector(to_unsigned(38, 8)),
			731 => std_logic_vector(to_unsigned(39, 8)),
			732 => std_logic_vector(to_unsigned(96, 8)),
			733 => std_logic_vector(to_unsigned(104, 8)),
			734 => std_logic_vector(to_unsigned(116, 8)),
			735 => std_logic_vector(to_unsigned(60, 8)),
			736 => std_logic_vector(to_unsigned(74, 8)),
			737 => std_logic_vector(to_unsigned(239, 8)),
			738 => std_logic_vector(to_unsigned(114, 8)),
			739 => std_logic_vector(to_unsigned(95, 8)),
			740 => std_logic_vector(to_unsigned(184, 8)),
			741 => std_logic_vector(to_unsigned(172, 8)),
			742 => std_logic_vector(to_unsigned(224, 8)),
			743 => std_logic_vector(to_unsigned(167, 8)),
			744 => std_logic_vector(to_unsigned(163, 8)),
			745 => std_logic_vector(to_unsigned(13, 8)),
			746 => std_logic_vector(to_unsigned(225, 8)),
			747 => std_logic_vector(to_unsigned(122, 8)),
			748 => std_logic_vector(to_unsigned(26, 8)),
			749 => std_logic_vector(to_unsigned(212, 8)),
			750 => std_logic_vector(to_unsigned(8, 8)),
			751 => std_logic_vector(to_unsigned(108, 8)),
			752 => std_logic_vector(to_unsigned(43, 8)),
			753 => std_logic_vector(to_unsigned(173, 8)),
			754 => std_logic_vector(to_unsigned(218, 8)),
			755 => std_logic_vector(to_unsigned(251, 8)),
			756 => std_logic_vector(to_unsigned(33, 8)),
			757 => std_logic_vector(to_unsigned(119, 8)),
			758 => std_logic_vector(to_unsigned(2, 8)),
			759 => std_logic_vector(to_unsigned(59, 8)),
			760 => std_logic_vector(to_unsigned(154, 8)),
			761 => std_logic_vector(to_unsigned(119, 8)),
			762 => std_logic_vector(to_unsigned(85, 8)),
			763 => std_logic_vector(to_unsigned(72, 8)),
			764 => std_logic_vector(to_unsigned(196, 8)),
			765 => std_logic_vector(to_unsigned(191, 8)),
			766 => std_logic_vector(to_unsigned(202, 8)),
			767 => std_logic_vector(to_unsigned(155, 8)),
			768 => std_logic_vector(to_unsigned(23, 8)),
			769 => std_logic_vector(to_unsigned(9, 8)),
			770 => std_logic_vector(to_unsigned(167, 8)),
			771 => std_logic_vector(to_unsigned(141, 8)),
			772 => std_logic_vector(to_unsigned(32, 8)),
			773 => std_logic_vector(to_unsigned(179, 8)),
			774 => std_logic_vector(to_unsigned(177, 8)),
			775 => std_logic_vector(to_unsigned(107, 8)),
			776 => std_logic_vector(to_unsigned(195, 8)),
			777 => std_logic_vector(to_unsigned(114, 8)),
			778 => std_logic_vector(to_unsigned(67, 8)),
			779 => std_logic_vector(to_unsigned(251, 8)),
			780 => std_logic_vector(to_unsigned(234, 8)),
			781 => std_logic_vector(to_unsigned(17, 8)),
			782 => std_logic_vector(to_unsigned(135, 8)),
			783 => std_logic_vector(to_unsigned(255, 8)),
			784 => std_logic_vector(to_unsigned(234, 8)),
			785 => std_logic_vector(to_unsigned(128, 8)),
			786 => std_logic_vector(to_unsigned(19, 8)),
			787 => std_logic_vector(to_unsigned(87, 8)),
			788 => std_logic_vector(to_unsigned(224, 8)),
			789 => std_logic_vector(to_unsigned(229, 8)),
			790 => std_logic_vector(to_unsigned(6, 8)),
			791 => std_logic_vector(to_unsigned(111, 8)),
			792 => std_logic_vector(to_unsigned(195, 8)),
			793 => std_logic_vector(to_unsigned(118, 8)),
			794 => std_logic_vector(to_unsigned(176, 8)),
			795 => std_logic_vector(to_unsigned(92, 8)),
			796 => std_logic_vector(to_unsigned(82, 8)),
			797 => std_logic_vector(to_unsigned(61, 8)),
			798 => std_logic_vector(to_unsigned(137, 8)),
			799 => std_logic_vector(to_unsigned(199, 8)),
			800 => std_logic_vector(to_unsigned(25, 8)),
			801 => std_logic_vector(to_unsigned(47, 8)),
			802 => std_logic_vector(to_unsigned(112, 8)),
			803 => std_logic_vector(to_unsigned(81, 8)),
			804 => std_logic_vector(to_unsigned(233, 8)),
			805 => std_logic_vector(to_unsigned(255, 8)),
			806 => std_logic_vector(to_unsigned(139, 8)),
			807 => std_logic_vector(to_unsigned(45, 8)),
			808 => std_logic_vector(to_unsigned(176, 8)),
			809 => std_logic_vector(to_unsigned(69, 8)),
			810 => std_logic_vector(to_unsigned(142, 8)),
			811 => std_logic_vector(to_unsigned(166, 8)),
			812 => std_logic_vector(to_unsigned(84, 8)),
			813 => std_logic_vector(to_unsigned(80, 8)),
			814 => std_logic_vector(to_unsigned(147, 8)),
			815 => std_logic_vector(to_unsigned(100, 8)),
			816 => std_logic_vector(to_unsigned(202, 8)),
			817 => std_logic_vector(to_unsigned(21, 8)),
			818 => std_logic_vector(to_unsigned(76, 8)),
			819 => std_logic_vector(to_unsigned(105, 8)),
			820 => std_logic_vector(to_unsigned(107, 8)),
			821 => std_logic_vector(to_unsigned(91, 8)),
			822 => std_logic_vector(to_unsigned(93, 8)),
			823 => std_logic_vector(to_unsigned(127, 8)),
			824 => std_logic_vector(to_unsigned(66, 8)),
			825 => std_logic_vector(to_unsigned(198, 8)),
			826 => std_logic_vector(to_unsigned(18, 8)),
			827 => std_logic_vector(to_unsigned(32, 8)),
			828 => std_logic_vector(to_unsigned(96, 8)),
			829 => std_logic_vector(to_unsigned(5, 8)),
			830 => std_logic_vector(to_unsigned(209, 8)),
			831 => std_logic_vector(to_unsigned(34, 8)),
			832 => std_logic_vector(to_unsigned(209, 8)),
			833 => std_logic_vector(to_unsigned(88, 8)),
			834 => std_logic_vector(to_unsigned(109, 8)),
			835 => std_logic_vector(to_unsigned(235, 8)),
			836 => std_logic_vector(to_unsigned(105, 8)),
			837 => std_logic_vector(to_unsigned(63, 8)),
			838 => std_logic_vector(to_unsigned(244, 8)),
			839 => std_logic_vector(to_unsigned(50, 8)),
			840 => std_logic_vector(to_unsigned(37, 8)),
			841 => std_logic_vector(to_unsigned(36, 8)),
			842 => std_logic_vector(to_unsigned(254, 8)),
			843 => std_logic_vector(to_unsigned(163, 8)),
			844 => std_logic_vector(to_unsigned(24, 8)),
			845 => std_logic_vector(to_unsigned(187, 8)),
			846 => std_logic_vector(to_unsigned(217, 8)),
			847 => std_logic_vector(to_unsigned(22, 8)),
			848 => std_logic_vector(to_unsigned(198, 8)),
			849 => std_logic_vector(to_unsigned(200, 8)),
			850 => std_logic_vector(to_unsigned(147, 8)),
			851 => std_logic_vector(to_unsigned(224, 8)),
			852 => std_logic_vector(to_unsigned(134, 8)),
			853 => std_logic_vector(to_unsigned(112, 8)),
			854 => std_logic_vector(to_unsigned(162, 8)),
			855 => std_logic_vector(to_unsigned(184, 8)),
			856 => std_logic_vector(to_unsigned(193, 8)),
			857 => std_logic_vector(to_unsigned(51, 8)),
			858 => std_logic_vector(to_unsigned(22, 8)),
			859 => std_logic_vector(to_unsigned(113, 8)),
			860 => std_logic_vector(to_unsigned(212, 8)),
			861 => std_logic_vector(to_unsigned(37, 8)),
			862 => std_logic_vector(to_unsigned(48, 8)),
			863 => std_logic_vector(to_unsigned(248, 8)),
			864 => std_logic_vector(to_unsigned(148, 8)),
			865 => std_logic_vector(to_unsigned(220, 8)),
			866 => std_logic_vector(to_unsigned(129, 8)),
			867 => std_logic_vector(to_unsigned(25, 8)),
			868 => std_logic_vector(to_unsigned(188, 8)),
			869 => std_logic_vector(to_unsigned(7, 8)),
			870 => std_logic_vector(to_unsigned(123, 8)),
			871 => std_logic_vector(to_unsigned(125, 8)),
			872 => std_logic_vector(to_unsigned(19, 8)),
			873 => std_logic_vector(to_unsigned(36, 8)),
			874 => std_logic_vector(to_unsigned(204, 8)),
			875 => std_logic_vector(to_unsigned(132, 8)),
			876 => std_logic_vector(to_unsigned(242, 8)),
			877 => std_logic_vector(to_unsigned(130, 8)),
			878 => std_logic_vector(to_unsigned(69, 8)),
			879 => std_logic_vector(to_unsigned(145, 8)),
			880 => std_logic_vector(to_unsigned(71, 8)),
			881 => std_logic_vector(to_unsigned(244, 8)),
			882 => std_logic_vector(to_unsigned(69, 8)),
			883 => std_logic_vector(to_unsigned(45, 8)),
			884 => std_logic_vector(to_unsigned(2, 8)),
			885 => std_logic_vector(to_unsigned(121, 8)),
			886 => std_logic_vector(to_unsigned(44, 8)),
			887 => std_logic_vector(to_unsigned(178, 8)),
			888 => std_logic_vector(to_unsigned(5, 8)),
			889 => std_logic_vector(to_unsigned(91, 8)),
			890 => std_logic_vector(to_unsigned(216, 8)),
			891 => std_logic_vector(to_unsigned(53, 8)),
			892 => std_logic_vector(to_unsigned(203, 8)),
			893 => std_logic_vector(to_unsigned(70, 8)),
			894 => std_logic_vector(to_unsigned(205, 8)),
			895 => std_logic_vector(to_unsigned(76, 8)),
			896 => std_logic_vector(to_unsigned(151, 8)),
			897 => std_logic_vector(to_unsigned(26, 8)),
			898 => std_logic_vector(to_unsigned(45, 8)),
			899 => std_logic_vector(to_unsigned(247, 8)),
			900 => std_logic_vector(to_unsigned(90, 8)),
			901 => std_logic_vector(to_unsigned(248, 8)),
			902 => std_logic_vector(to_unsigned(34, 8)),
			903 => std_logic_vector(to_unsigned(203, 8)),
			904 => std_logic_vector(to_unsigned(79, 8)),
			905 => std_logic_vector(to_unsigned(193, 8)),
			906 => std_logic_vector(to_unsigned(235, 8)),
			907 => std_logic_vector(to_unsigned(89, 8)),
			908 => std_logic_vector(to_unsigned(205, 8)),
			909 => std_logic_vector(to_unsigned(227, 8)),
			910 => std_logic_vector(to_unsigned(26, 8)),
			911 => std_logic_vector(to_unsigned(133, 8)),
			912 => std_logic_vector(to_unsigned(95, 8)),
			913 => std_logic_vector(to_unsigned(203, 8)),
			914 => std_logic_vector(to_unsigned(89, 8)),
			915 => std_logic_vector(to_unsigned(165, 8)),
			916 => std_logic_vector(to_unsigned(244, 8)),
			917 => std_logic_vector(to_unsigned(132, 8)),
			918 => std_logic_vector(to_unsigned(82, 8)),
			919 => std_logic_vector(to_unsigned(200, 8)),
			920 => std_logic_vector(to_unsigned(237, 8)),
			921 => std_logic_vector(to_unsigned(98, 8)),
			922 => std_logic_vector(to_unsigned(222, 8)),
			923 => std_logic_vector(to_unsigned(8, 8)),
			924 => std_logic_vector(to_unsigned(239, 8)),
			925 => std_logic_vector(to_unsigned(112, 8)),
			926 => std_logic_vector(to_unsigned(158, 8)),
			927 => std_logic_vector(to_unsigned(151, 8)),
			928 => std_logic_vector(to_unsigned(51, 8)),
			929 => std_logic_vector(to_unsigned(248, 8)),
			930 => std_logic_vector(to_unsigned(210, 8)),
			931 => std_logic_vector(to_unsigned(20, 8)),
			932 => std_logic_vector(to_unsigned(15, 8)),
			933 => std_logic_vector(to_unsigned(160, 8)),
			934 => std_logic_vector(to_unsigned(92, 8)),
			935 => std_logic_vector(to_unsigned(36, 8)),
			936 => std_logic_vector(to_unsigned(39, 8)),
			937 => std_logic_vector(to_unsigned(155, 8)),
			938 => std_logic_vector(to_unsigned(50, 8)),
			939 => std_logic_vector(to_unsigned(145, 8)),
			940 => std_logic_vector(to_unsigned(224, 8)),
			941 => std_logic_vector(to_unsigned(250, 8)),
			942 => std_logic_vector(to_unsigned(242, 8)),
			943 => std_logic_vector(to_unsigned(109, 8)),
			944 => std_logic_vector(to_unsigned(44, 8)),
			945 => std_logic_vector(to_unsigned(26, 8)),
			946 => std_logic_vector(to_unsigned(112, 8)),
			947 => std_logic_vector(to_unsigned(106, 8)),
			948 => std_logic_vector(to_unsigned(200, 8)),
			949 => std_logic_vector(to_unsigned(46, 8)),
			950 => std_logic_vector(to_unsigned(170, 8)),
			951 => std_logic_vector(to_unsigned(72, 8)),
			952 => std_logic_vector(to_unsigned(100, 8)),
			953 => std_logic_vector(to_unsigned(23, 8)),
			954 => std_logic_vector(to_unsigned(217, 8)),
			955 => std_logic_vector(to_unsigned(222, 8)),
			956 => std_logic_vector(to_unsigned(20, 8)),
			957 => std_logic_vector(to_unsigned(105, 8)),
			958 => std_logic_vector(to_unsigned(255, 8)),
			959 => std_logic_vector(to_unsigned(181, 8)),
			960 => std_logic_vector(to_unsigned(233, 8)),
			961 => std_logic_vector(to_unsigned(35, 8)),
			962 => std_logic_vector(to_unsigned(207, 8)),
			963 => std_logic_vector(to_unsigned(24, 8)),
			964 => std_logic_vector(to_unsigned(222, 8)),
			965 => std_logic_vector(to_unsigned(92, 8)),
			966 => std_logic_vector(to_unsigned(172, 8)),
			967 => std_logic_vector(to_unsigned(24, 8)),
			968 => std_logic_vector(to_unsigned(85, 8)),
			969 => std_logic_vector(to_unsigned(29, 8)),
			970 => std_logic_vector(to_unsigned(80, 8)),
			971 => std_logic_vector(to_unsigned(67, 8)),
			972 => std_logic_vector(to_unsigned(47, 8)),
			973 => std_logic_vector(to_unsigned(184, 8)),
			974 => std_logic_vector(to_unsigned(193, 8)),
			975 => std_logic_vector(to_unsigned(254, 8)),
			976 => std_logic_vector(to_unsigned(137, 8)),
			977 => std_logic_vector(to_unsigned(145, 8)),
			978 => std_logic_vector(to_unsigned(97, 8)),
			979 => std_logic_vector(to_unsigned(232, 8)),
			980 => std_logic_vector(to_unsigned(220, 8)),
			981 => std_logic_vector(to_unsigned(75, 8)),
			982 => std_logic_vector(to_unsigned(88, 8)),
			983 => std_logic_vector(to_unsigned(56, 8)),
			984 => std_logic_vector(to_unsigned(226, 8)),
			985 => std_logic_vector(to_unsigned(234, 8)),
			986 => std_logic_vector(to_unsigned(56, 8)),
			987 => std_logic_vector(to_unsigned(158, 8)),
			988 => std_logic_vector(to_unsigned(27, 8)),
			989 => std_logic_vector(to_unsigned(104, 8)),
			990 => std_logic_vector(to_unsigned(169, 8)),
			991 => std_logic_vector(to_unsigned(134, 8)),
			992 => std_logic_vector(to_unsigned(7, 8)),
			993 => std_logic_vector(to_unsigned(160, 8)),
			994 => std_logic_vector(to_unsigned(182, 8)),
			995 => std_logic_vector(to_unsigned(32, 8)),
			996 => std_logic_vector(to_unsigned(44, 8)),
			997 => std_logic_vector(to_unsigned(127, 8)),
			998 => std_logic_vector(to_unsigned(193, 8)),
			999 => std_logic_vector(to_unsigned(101, 8)),
			1000 => std_logic_vector(to_unsigned(205, 8)),
			1001 => std_logic_vector(to_unsigned(2, 8)),
			1002 => std_logic_vector(to_unsigned(200, 8)),
			1003 => std_logic_vector(to_unsigned(194, 8)),
			1004 => std_logic_vector(to_unsigned(184, 8)),
			1005 => std_logic_vector(to_unsigned(96, 8)),
			1006 => std_logic_vector(to_unsigned(96, 8)),
			1007 => std_logic_vector(to_unsigned(221, 8)),
			1008 => std_logic_vector(to_unsigned(18, 8)),
			1009 => std_logic_vector(to_unsigned(102, 8)),
			1010 => std_logic_vector(to_unsigned(24, 8)),
			1011 => std_logic_vector(to_unsigned(148, 8)),
			1012 => std_logic_vector(to_unsigned(99, 8)),
			1013 => std_logic_vector(to_unsigned(32, 8)),
			1014 => std_logic_vector(to_unsigned(227, 8)),
			1015 => std_logic_vector(to_unsigned(65, 8)),
			1016 => std_logic_vector(to_unsigned(164, 8)),
			1017 => std_logic_vector(to_unsigned(97, 8)),
			1018 => std_logic_vector(to_unsigned(14, 8)),
			1019 => std_logic_vector(to_unsigned(183, 8)),
			1020 => std_logic_vector(to_unsigned(13, 8)),
			1021 => std_logic_vector(to_unsigned(186, 8)),
			1022 => std_logic_vector(to_unsigned(229, 8)),
			1023 => std_logic_vector(to_unsigned(192, 8)),
			1024 => std_logic_vector(to_unsigned(115, 8)),
			1025 => std_logic_vector(to_unsigned(157, 8)),
			1026 => std_logic_vector(to_unsigned(218, 8)),
			1027 => std_logic_vector(to_unsigned(236, 8)),
			1028 => std_logic_vector(to_unsigned(124, 8)),
			1029 => std_logic_vector(to_unsigned(173, 8)),
			1030 => std_logic_vector(to_unsigned(138, 8)),
			1031 => std_logic_vector(to_unsigned(230, 8)),
			1032 => std_logic_vector(to_unsigned(47, 8)),
			1033 => std_logic_vector(to_unsigned(201, 8)),
			1034 => std_logic_vector(to_unsigned(126, 8)),
			1035 => std_logic_vector(to_unsigned(117, 8)),
			1036 => std_logic_vector(to_unsigned(127, 8)),
			1037 => std_logic_vector(to_unsigned(243, 8)),
			1038 => std_logic_vector(to_unsigned(6, 8)),
			1039 => std_logic_vector(to_unsigned(110, 8)),
			1040 => std_logic_vector(to_unsigned(93, 8)),
			1041 => std_logic_vector(to_unsigned(84, 8)),
			1042 => std_logic_vector(to_unsigned(98, 8)),
			1043 => std_logic_vector(to_unsigned(125, 8)),
			1044 => std_logic_vector(to_unsigned(214, 8)),
			1045 => std_logic_vector(to_unsigned(111, 8)),
			1046 => std_logic_vector(to_unsigned(176, 8)),
			1047 => std_logic_vector(to_unsigned(190, 8)),
			1048 => std_logic_vector(to_unsigned(106, 8)),
			1049 => std_logic_vector(to_unsigned(42, 8)),
			1050 => std_logic_vector(to_unsigned(217, 8)),
			1051 => std_logic_vector(to_unsigned(185, 8)),
			1052 => std_logic_vector(to_unsigned(37, 8)),
			1053 => std_logic_vector(to_unsigned(85, 8)),
			1054 => std_logic_vector(to_unsigned(50, 8)),
			1055 => std_logic_vector(to_unsigned(72, 8)),
			1056 => std_logic_vector(to_unsigned(89, 8)),
			1057 => std_logic_vector(to_unsigned(23, 8)),
			1058 => std_logic_vector(to_unsigned(143, 8)),
			1059 => std_logic_vector(to_unsigned(195, 8)),
			1060 => std_logic_vector(to_unsigned(249, 8)),
			1061 => std_logic_vector(to_unsigned(87, 8)),
			1062 => std_logic_vector(to_unsigned(81, 8)),
			1063 => std_logic_vector(to_unsigned(199, 8)),
			1064 => std_logic_vector(to_unsigned(120, 8)),
			1065 => std_logic_vector(to_unsigned(85, 8)),
			1066 => std_logic_vector(to_unsigned(121, 8)),
			1067 => std_logic_vector(to_unsigned(17, 8)),
			1068 => std_logic_vector(to_unsigned(225, 8)),
			1069 => std_logic_vector(to_unsigned(195, 8)),
			1070 => std_logic_vector(to_unsigned(177, 8)),
			1071 => std_logic_vector(to_unsigned(196, 8)),
			1072 => std_logic_vector(to_unsigned(81, 8)),
			1073 => std_logic_vector(to_unsigned(192, 8)),
			1074 => std_logic_vector(to_unsigned(253, 8)),
			1075 => std_logic_vector(to_unsigned(59, 8)),
			1076 => std_logic_vector(to_unsigned(113, 8)),
			1077 => std_logic_vector(to_unsigned(44, 8)),
			1078 => std_logic_vector(to_unsigned(98, 8)),
			1079 => std_logic_vector(to_unsigned(54, 8)),
			1080 => std_logic_vector(to_unsigned(223, 8)),
			1081 => std_logic_vector(to_unsigned(50, 8)),
			1082 => std_logic_vector(to_unsigned(49, 8)),
			1083 => std_logic_vector(to_unsigned(135, 8)),
			1084 => std_logic_vector(to_unsigned(80, 8)),
			1085 => std_logic_vector(to_unsigned(48, 8)),
			1086 => std_logic_vector(to_unsigned(233, 8)),
			1087 => std_logic_vector(to_unsigned(21, 8)),
			1088 => std_logic_vector(to_unsigned(134, 8)),
			1089 => std_logic_vector(to_unsigned(49, 8)),
			1090 => std_logic_vector(to_unsigned(254, 8)),
			1091 => std_logic_vector(to_unsigned(177, 8)),
			1092 => std_logic_vector(to_unsigned(146, 8)),
			1093 => std_logic_vector(to_unsigned(50, 8)),
			1094 => std_logic_vector(to_unsigned(135, 8)),
			1095 => std_logic_vector(to_unsigned(117, 8)),
			1096 => std_logic_vector(to_unsigned(222, 8)),
			1097 => std_logic_vector(to_unsigned(174, 8)),
			1098 => std_logic_vector(to_unsigned(238, 8)),
			1099 => std_logic_vector(to_unsigned(248, 8)),
			1100 => std_logic_vector(to_unsigned(193, 8)),
			1101 => std_logic_vector(to_unsigned(193, 8)),
			1102 => std_logic_vector(to_unsigned(203, 8)),
			1103 => std_logic_vector(to_unsigned(200, 8)),
			1104 => std_logic_vector(to_unsigned(102, 8)),
			1105 => std_logic_vector(to_unsigned(186, 8)),
			1106 => std_logic_vector(to_unsigned(6, 8)),
			1107 => std_logic_vector(to_unsigned(122, 8)),
			1108 => std_logic_vector(to_unsigned(82, 8)),
			1109 => std_logic_vector(to_unsigned(125, 8)),
			1110 => std_logic_vector(to_unsigned(19, 8)),
			1111 => std_logic_vector(to_unsigned(125, 8)),
			1112 => std_logic_vector(to_unsigned(248, 8)),
			1113 => std_logic_vector(to_unsigned(134, 8)),
			1114 => std_logic_vector(to_unsigned(174, 8)),
			1115 => std_logic_vector(to_unsigned(182, 8)),
			1116 => std_logic_vector(to_unsigned(33, 8)),
			1117 => std_logic_vector(to_unsigned(235, 8)),
			1118 => std_logic_vector(to_unsigned(36, 8)),
			1119 => std_logic_vector(to_unsigned(146, 8)),
			1120 => std_logic_vector(to_unsigned(5, 8)),
			1121 => std_logic_vector(to_unsigned(205, 8)),
			1122 => std_logic_vector(to_unsigned(243, 8)),
			1123 => std_logic_vector(to_unsigned(184, 8)),
			1124 => std_logic_vector(to_unsigned(148, 8)),
			1125 => std_logic_vector(to_unsigned(81, 8)),
			1126 => std_logic_vector(to_unsigned(211, 8)),
			1127 => std_logic_vector(to_unsigned(195, 8)),
			1128 => std_logic_vector(to_unsigned(72, 8)),
			1129 => std_logic_vector(to_unsigned(221, 8)),
			1130 => std_logic_vector(to_unsigned(142, 8)),
			1131 => std_logic_vector(to_unsigned(182, 8)),
			1132 => std_logic_vector(to_unsigned(7, 8)),
			1133 => std_logic_vector(to_unsigned(237, 8)),
			1134 => std_logic_vector(to_unsigned(62, 8)),
			1135 => std_logic_vector(to_unsigned(223, 8)),
			1136 => std_logic_vector(to_unsigned(61, 8)),
			1137 => std_logic_vector(to_unsigned(135, 8)),
			1138 => std_logic_vector(to_unsigned(66, 8)),
			1139 => std_logic_vector(to_unsigned(123, 8)),
			1140 => std_logic_vector(to_unsigned(202, 8)),
			1141 => std_logic_vector(to_unsigned(46, 8)),
			1142 => std_logic_vector(to_unsigned(171, 8)),
			1143 => std_logic_vector(to_unsigned(34, 8)),
			1144 => std_logic_vector(to_unsigned(35, 8)),
			1145 => std_logic_vector(to_unsigned(167, 8)),
			1146 => std_logic_vector(to_unsigned(75, 8)),
			1147 => std_logic_vector(to_unsigned(91, 8)),
			1148 => std_logic_vector(to_unsigned(49, 8)),
			1149 => std_logic_vector(to_unsigned(36, 8)),
			1150 => std_logic_vector(to_unsigned(101, 8)),
			1151 => std_logic_vector(to_unsigned(50, 8)),
			1152 => std_logic_vector(to_unsigned(209, 8)),
			1153 => std_logic_vector(to_unsigned(215, 8)),
			1154 => std_logic_vector(to_unsigned(147, 8)),
			1155 => std_logic_vector(to_unsigned(78, 8)),
			1156 => std_logic_vector(to_unsigned(224, 8)),
			1157 => std_logic_vector(to_unsigned(205, 8)),
			1158 => std_logic_vector(to_unsigned(251, 8)),
			1159 => std_logic_vector(to_unsigned(186, 8)),
			1160 => std_logic_vector(to_unsigned(151, 8)),
			1161 => std_logic_vector(to_unsigned(219, 8)),
			1162 => std_logic_vector(to_unsigned(230, 8)),
			1163 => std_logic_vector(to_unsigned(213, 8)),
			1164 => std_logic_vector(to_unsigned(181, 8)),
			1165 => std_logic_vector(to_unsigned(188, 8)),
			1166 => std_logic_vector(to_unsigned(224, 8)),
			1167 => std_logic_vector(to_unsigned(89, 8)),
			1168 => std_logic_vector(to_unsigned(213, 8)),
			1169 => std_logic_vector(to_unsigned(143, 8)),
			1170 => std_logic_vector(to_unsigned(201, 8)),
			1171 => std_logic_vector(to_unsigned(113, 8)),
			1172 => std_logic_vector(to_unsigned(47, 8)),
			1173 => std_logic_vector(to_unsigned(191, 8)),
			1174 => std_logic_vector(to_unsigned(223, 8)),
			1175 => std_logic_vector(to_unsigned(199, 8)),
			1176 => std_logic_vector(to_unsigned(218, 8)),
			1177 => std_logic_vector(to_unsigned(108, 8)),
			1178 => std_logic_vector(to_unsigned(31, 8)),
			1179 => std_logic_vector(to_unsigned(38, 8)),
			1180 => std_logic_vector(to_unsigned(63, 8)),
			1181 => std_logic_vector(to_unsigned(174, 8)),
			1182 => std_logic_vector(to_unsigned(11, 8)),
			1183 => std_logic_vector(to_unsigned(25, 8)),
			1184 => std_logic_vector(to_unsigned(93, 8)),
			1185 => std_logic_vector(to_unsigned(236, 8)),
			1186 => std_logic_vector(to_unsigned(182, 8)),
			1187 => std_logic_vector(to_unsigned(163, 8)),
			1188 => std_logic_vector(to_unsigned(110, 8)),
			1189 => std_logic_vector(to_unsigned(10, 8)),
			1190 => std_logic_vector(to_unsigned(43, 8)),
			1191 => std_logic_vector(to_unsigned(118, 8)),
			1192 => std_logic_vector(to_unsigned(102, 8)),
			1193 => std_logic_vector(to_unsigned(158, 8)),
			1194 => std_logic_vector(to_unsigned(78, 8)),
			1195 => std_logic_vector(to_unsigned(228, 8)),
			1196 => std_logic_vector(to_unsigned(177, 8)),
			1197 => std_logic_vector(to_unsigned(137, 8)),
			1198 => std_logic_vector(to_unsigned(36, 8)),
			1199 => std_logic_vector(to_unsigned(200, 8)),
			1200 => std_logic_vector(to_unsigned(78, 8)),
			1201 => std_logic_vector(to_unsigned(152, 8)),
			1202 => std_logic_vector(to_unsigned(61, 8)),
			1203 => std_logic_vector(to_unsigned(153, 8)),
			1204 => std_logic_vector(to_unsigned(150, 8)),
			1205 => std_logic_vector(to_unsigned(76, 8)),
			1206 => std_logic_vector(to_unsigned(62, 8)),
			1207 => std_logic_vector(to_unsigned(165, 8)),
			1208 => std_logic_vector(to_unsigned(57, 8)),
			1209 => std_logic_vector(to_unsigned(178, 8)),
			1210 => std_logic_vector(to_unsigned(254, 8)),
			1211 => std_logic_vector(to_unsigned(183, 8)),
			1212 => std_logic_vector(to_unsigned(70, 8)),
			1213 => std_logic_vector(to_unsigned(120, 8)),
			1214 => std_logic_vector(to_unsigned(39, 8)),
			1215 => std_logic_vector(to_unsigned(38, 8)),
			1216 => std_logic_vector(to_unsigned(141, 8)),
			1217 => std_logic_vector(to_unsigned(60, 8)),
			1218 => std_logic_vector(to_unsigned(234, 8)),
			1219 => std_logic_vector(to_unsigned(157, 8)),
			1220 => std_logic_vector(to_unsigned(223, 8)),
			1221 => std_logic_vector(to_unsigned(184, 8)),
			1222 => std_logic_vector(to_unsigned(35, 8)),
			1223 => std_logic_vector(to_unsigned(252, 8)),
			1224 => std_logic_vector(to_unsigned(155, 8)),
			1225 => std_logic_vector(to_unsigned(252, 8)),
			1226 => std_logic_vector(to_unsigned(143, 8)),
			1227 => std_logic_vector(to_unsigned(201, 8)),
			1228 => std_logic_vector(to_unsigned(174, 8)),
			1229 => std_logic_vector(to_unsigned(51, 8)),
			1230 => std_logic_vector(to_unsigned(12, 8)),
			1231 => std_logic_vector(to_unsigned(223, 8)),
			1232 => std_logic_vector(to_unsigned(5, 8)),
			1233 => std_logic_vector(to_unsigned(102, 8)),
			1234 => std_logic_vector(to_unsigned(67, 8)),
			1235 => std_logic_vector(to_unsigned(249, 8)),
			1236 => std_logic_vector(to_unsigned(146, 8)),
			1237 => std_logic_vector(to_unsigned(30, 8)),
			1238 => std_logic_vector(to_unsigned(177, 8)),
			1239 => std_logic_vector(to_unsigned(76, 8)),
			1240 => std_logic_vector(to_unsigned(218, 8)),
			1241 => std_logic_vector(to_unsigned(149, 8)),
			1242 => std_logic_vector(to_unsigned(69, 8)),
			1243 => std_logic_vector(to_unsigned(84, 8)),
			1244 => std_logic_vector(to_unsigned(141, 8)),
			1245 => std_logic_vector(to_unsigned(13, 8)),
			1246 => std_logic_vector(to_unsigned(152, 8)),
			1247 => std_logic_vector(to_unsigned(143, 8)),
			1248 => std_logic_vector(to_unsigned(246, 8)),
			1249 => std_logic_vector(to_unsigned(125, 8)),
			1250 => std_logic_vector(to_unsigned(73, 8)),
			1251 => std_logic_vector(to_unsigned(108, 8)),
			1252 => std_logic_vector(to_unsigned(88, 8)),
			1253 => std_logic_vector(to_unsigned(10, 8)),
			1254 => std_logic_vector(to_unsigned(241, 8)),
			1255 => std_logic_vector(to_unsigned(248, 8)),
			1256 => std_logic_vector(to_unsigned(251, 8)),
			1257 => std_logic_vector(to_unsigned(183, 8)),
			1258 => std_logic_vector(to_unsigned(123, 8)),
			1259 => std_logic_vector(to_unsigned(94, 8)),
			1260 => std_logic_vector(to_unsigned(64, 8)),
			1261 => std_logic_vector(to_unsigned(244, 8)),
			1262 => std_logic_vector(to_unsigned(216, 8)),
			1263 => std_logic_vector(to_unsigned(241, 8)),
			1264 => std_logic_vector(to_unsigned(9, 8)),
			1265 => std_logic_vector(to_unsigned(117, 8)),
			1266 => std_logic_vector(to_unsigned(213, 8)),
			1267 => std_logic_vector(to_unsigned(105, 8)),
			1268 => std_logic_vector(to_unsigned(183, 8)),
			1269 => std_logic_vector(to_unsigned(52, 8)),
			1270 => std_logic_vector(to_unsigned(95, 8)),
			1271 => std_logic_vector(to_unsigned(210, 8)),
			1272 => std_logic_vector(to_unsigned(245, 8)),
			1273 => std_logic_vector(to_unsigned(27, 8)),
			1274 => std_logic_vector(to_unsigned(27, 8)),
			1275 => std_logic_vector(to_unsigned(20, 8)),
			1276 => std_logic_vector(to_unsigned(46, 8)),
			1277 => std_logic_vector(to_unsigned(151, 8)),
			1278 => std_logic_vector(to_unsigned(121, 8)),
			1279 => std_logic_vector(to_unsigned(141, 8)),
			1280 => std_logic_vector(to_unsigned(193, 8)),
			1281 => std_logic_vector(to_unsigned(47, 8)),
			1282 => std_logic_vector(to_unsigned(218, 8)),
			1283 => std_logic_vector(to_unsigned(117, 8)),
			1284 => std_logic_vector(to_unsigned(23, 8)),
			1285 => std_logic_vector(to_unsigned(56, 8)),
			1286 => std_logic_vector(to_unsigned(178, 8)),
			1287 => std_logic_vector(to_unsigned(155, 8)),
			1288 => std_logic_vector(to_unsigned(240, 8)),
			1289 => std_logic_vector(to_unsigned(135, 8)),
			1290 => std_logic_vector(to_unsigned(119, 8)),
			1291 => std_logic_vector(to_unsigned(72, 8)),
			1292 => std_logic_vector(to_unsigned(90, 8)),
			1293 => std_logic_vector(to_unsigned(72, 8)),
			1294 => std_logic_vector(to_unsigned(26, 8)),
			1295 => std_logic_vector(to_unsigned(16, 8)),
			1296 => std_logic_vector(to_unsigned(110, 8)),
			1297 => std_logic_vector(to_unsigned(228, 8)),
			1298 => std_logic_vector(to_unsigned(178, 8)),
			1299 => std_logic_vector(to_unsigned(20, 8)),
			1300 => std_logic_vector(to_unsigned(121, 8)),
			1301 => std_logic_vector(to_unsigned(163, 8)),
			1302 => std_logic_vector(to_unsigned(154, 8)),
			1303 => std_logic_vector(to_unsigned(66, 8)),
			1304 => std_logic_vector(to_unsigned(181, 8)),
			1305 => std_logic_vector(to_unsigned(90, 8)),
			1306 => std_logic_vector(to_unsigned(19, 8)),
			1307 => std_logic_vector(to_unsigned(73, 8)),
			1308 => std_logic_vector(to_unsigned(37, 8)),
			1309 => std_logic_vector(to_unsigned(29, 8)),
			1310 => std_logic_vector(to_unsigned(60, 8)),
			1311 => std_logic_vector(to_unsigned(237, 8)),
			1312 => std_logic_vector(to_unsigned(235, 8)),
			1313 => std_logic_vector(to_unsigned(30, 8)),
			1314 => std_logic_vector(to_unsigned(38, 8)),
			1315 => std_logic_vector(to_unsigned(216, 8)),
			1316 => std_logic_vector(to_unsigned(98, 8)),
			1317 => std_logic_vector(to_unsigned(82, 8)),
			1318 => std_logic_vector(to_unsigned(171, 8)),
			1319 => std_logic_vector(to_unsigned(158, 8)),
			1320 => std_logic_vector(to_unsigned(166, 8)),
			1321 => std_logic_vector(to_unsigned(183, 8)),
			1322 => std_logic_vector(to_unsigned(72, 8)),
			1323 => std_logic_vector(to_unsigned(76, 8)),
			1324 => std_logic_vector(to_unsigned(63, 8)),
			1325 => std_logic_vector(to_unsigned(99, 8)),
			1326 => std_logic_vector(to_unsigned(128, 8)),
			1327 => std_logic_vector(to_unsigned(144, 8)),
			1328 => std_logic_vector(to_unsigned(10, 8)),
			1329 => std_logic_vector(to_unsigned(101, 8)),
			1330 => std_logic_vector(to_unsigned(106, 8)),
			1331 => std_logic_vector(to_unsigned(160, 8)),
			1332 => std_logic_vector(to_unsigned(179, 8)),
			1333 => std_logic_vector(to_unsigned(90, 8)),
			1334 => std_logic_vector(to_unsigned(225, 8)),
			1335 => std_logic_vector(to_unsigned(109, 8)),
			1336 => std_logic_vector(to_unsigned(160, 8)),
			1337 => std_logic_vector(to_unsigned(117, 8)),
			1338 => std_logic_vector(to_unsigned(160, 8)),
			1339 => std_logic_vector(to_unsigned(245, 8)),
			1340 => std_logic_vector(to_unsigned(95, 8)),
			1341 => std_logic_vector(to_unsigned(14, 8)),
			1342 => std_logic_vector(to_unsigned(205, 8)),
			1343 => std_logic_vector(to_unsigned(144, 8)),
			1344 => std_logic_vector(to_unsigned(178, 8)),
			1345 => std_logic_vector(to_unsigned(3, 8)),
			1346 => std_logic_vector(to_unsigned(61, 8)),
			1347 => std_logic_vector(to_unsigned(127, 8)),
			1348 => std_logic_vector(to_unsigned(33, 8)),
			1349 => std_logic_vector(to_unsigned(3, 8)),
			1350 => std_logic_vector(to_unsigned(238, 8)),
			1351 => std_logic_vector(to_unsigned(96, 8)),
			1352 => std_logic_vector(to_unsigned(19, 8)),
			1353 => std_logic_vector(to_unsigned(191, 8)),
			1354 => std_logic_vector(to_unsigned(92, 8)),
			1355 => std_logic_vector(to_unsigned(156, 8)),
			1356 => std_logic_vector(to_unsigned(88, 8)),
			1357 => std_logic_vector(to_unsigned(134, 8)),
			1358 => std_logic_vector(to_unsigned(109, 8)),
			1359 => std_logic_vector(to_unsigned(23, 8)),
			1360 => std_logic_vector(to_unsigned(76, 8)),
			1361 => std_logic_vector(to_unsigned(241, 8)),
			1362 => std_logic_vector(to_unsigned(167, 8)),
			1363 => std_logic_vector(to_unsigned(215, 8)),
			1364 => std_logic_vector(to_unsigned(34, 8)),
			1365 => std_logic_vector(to_unsigned(143, 8)),
			1366 => std_logic_vector(to_unsigned(240, 8)),
			1367 => std_logic_vector(to_unsigned(78, 8)),
			1368 => std_logic_vector(to_unsigned(165, 8)),
			1369 => std_logic_vector(to_unsigned(178, 8)),
			1370 => std_logic_vector(to_unsigned(106, 8)),
			1371 => std_logic_vector(to_unsigned(12, 8)),
			1372 => std_logic_vector(to_unsigned(197, 8)),
			1373 => std_logic_vector(to_unsigned(32, 8)),
			1374 => std_logic_vector(to_unsigned(86, 8)),
			1375 => std_logic_vector(to_unsigned(61, 8)),
			1376 => std_logic_vector(to_unsigned(175, 8)),
			1377 => std_logic_vector(to_unsigned(90, 8)),
			1378 => std_logic_vector(to_unsigned(20, 8)),
			1379 => std_logic_vector(to_unsigned(117, 8)),
			1380 => std_logic_vector(to_unsigned(168, 8)),
			1381 => std_logic_vector(to_unsigned(118, 8)),
			1382 => std_logic_vector(to_unsigned(76, 8)),
			1383 => std_logic_vector(to_unsigned(38, 8)),
			1384 => std_logic_vector(to_unsigned(249, 8)),
			1385 => std_logic_vector(to_unsigned(250, 8)),
			1386 => std_logic_vector(to_unsigned(20, 8)),
			1387 => std_logic_vector(to_unsigned(20, 8)),
			1388 => std_logic_vector(to_unsigned(5, 8)),
			1389 => std_logic_vector(to_unsigned(192, 8)),
			1390 => std_logic_vector(to_unsigned(71, 8)),
			1391 => std_logic_vector(to_unsigned(131, 8)),
			1392 => std_logic_vector(to_unsigned(59, 8)),
			1393 => std_logic_vector(to_unsigned(53, 8)),
			1394 => std_logic_vector(to_unsigned(216, 8)),
			1395 => std_logic_vector(to_unsigned(141, 8)),
			1396 => std_logic_vector(to_unsigned(16, 8)),
			1397 => std_logic_vector(to_unsigned(149, 8)),
			1398 => std_logic_vector(to_unsigned(156, 8)),
			1399 => std_logic_vector(to_unsigned(108, 8)),
			1400 => std_logic_vector(to_unsigned(33, 8)),
			1401 => std_logic_vector(to_unsigned(150, 8)),
			1402 => std_logic_vector(to_unsigned(231, 8)),
			1403 => std_logic_vector(to_unsigned(156, 8)),
			1404 => std_logic_vector(to_unsigned(71, 8)),
			1405 => std_logic_vector(to_unsigned(216, 8)),
			1406 => std_logic_vector(to_unsigned(174, 8)),
			1407 => std_logic_vector(to_unsigned(109, 8)),
			1408 => std_logic_vector(to_unsigned(74, 8)),
			1409 => std_logic_vector(to_unsigned(158, 8)),
			1410 => std_logic_vector(to_unsigned(246, 8)),
			1411 => std_logic_vector(to_unsigned(116, 8)),
			1412 => std_logic_vector(to_unsigned(58, 8)),
			1413 => std_logic_vector(to_unsigned(113, 8)),
			1414 => std_logic_vector(to_unsigned(19, 8)),
			1415 => std_logic_vector(to_unsigned(183, 8)),
			1416 => std_logic_vector(to_unsigned(127, 8)),
			1417 => std_logic_vector(to_unsigned(247, 8)),
			1418 => std_logic_vector(to_unsigned(167, 8)),
			1419 => std_logic_vector(to_unsigned(214, 8)),
			1420 => std_logic_vector(to_unsigned(206, 8)),
			1421 => std_logic_vector(to_unsigned(243, 8)),
			1422 => std_logic_vector(to_unsigned(98, 8)),
			1423 => std_logic_vector(to_unsigned(246, 8)),
			1424 => std_logic_vector(to_unsigned(206, 8)),
			1425 => std_logic_vector(to_unsigned(252, 8)),
			1426 => std_logic_vector(to_unsigned(95, 8)),
			1427 => std_logic_vector(to_unsigned(128, 8)),
			1428 => std_logic_vector(to_unsigned(145, 8)),
			1429 => std_logic_vector(to_unsigned(24, 8)),
			1430 => std_logic_vector(to_unsigned(180, 8)),
			1431 => std_logic_vector(to_unsigned(166, 8)),
			1432 => std_logic_vector(to_unsigned(216, 8)),
			1433 => std_logic_vector(to_unsigned(126, 8)),
			1434 => std_logic_vector(to_unsigned(135, 8)),
			1435 => std_logic_vector(to_unsigned(57, 8)),
			1436 => std_logic_vector(to_unsigned(244, 8)),
			1437 => std_logic_vector(to_unsigned(132, 8)),
			1438 => std_logic_vector(to_unsigned(169, 8)),
			1439 => std_logic_vector(to_unsigned(104, 8)),
			1440 => std_logic_vector(to_unsigned(184, 8)),
			1441 => std_logic_vector(to_unsigned(154, 8)),
			1442 => std_logic_vector(to_unsigned(233, 8)),
			1443 => std_logic_vector(to_unsigned(74, 8)),
			1444 => std_logic_vector(to_unsigned(41, 8)),
			1445 => std_logic_vector(to_unsigned(254, 8)),
			1446 => std_logic_vector(to_unsigned(66, 8)),
			1447 => std_logic_vector(to_unsigned(32, 8)),
			1448 => std_logic_vector(to_unsigned(153, 8)),
			1449 => std_logic_vector(to_unsigned(78, 8)),
			1450 => std_logic_vector(to_unsigned(160, 8)),
			1451 => std_logic_vector(to_unsigned(212, 8)),
			1452 => std_logic_vector(to_unsigned(115, 8)),
			1453 => std_logic_vector(to_unsigned(34, 8)),
			1454 => std_logic_vector(to_unsigned(242, 8)),
			1455 => std_logic_vector(to_unsigned(46, 8)),
			1456 => std_logic_vector(to_unsigned(26, 8)),
			1457 => std_logic_vector(to_unsigned(110, 8)),
			1458 => std_logic_vector(to_unsigned(255, 8)),
			1459 => std_logic_vector(to_unsigned(48, 8)),
			1460 => std_logic_vector(to_unsigned(199, 8)),
			1461 => std_logic_vector(to_unsigned(42, 8)),
			1462 => std_logic_vector(to_unsigned(69, 8)),
			1463 => std_logic_vector(to_unsigned(57, 8)),
			1464 => std_logic_vector(to_unsigned(151, 8)),
			1465 => std_logic_vector(to_unsigned(206, 8)),
			1466 => std_logic_vector(to_unsigned(97, 8)),
			1467 => std_logic_vector(to_unsigned(189, 8)),
			1468 => std_logic_vector(to_unsigned(235, 8)),
			1469 => std_logic_vector(to_unsigned(217, 8)),
			1470 => std_logic_vector(to_unsigned(119, 8)),
			1471 => std_logic_vector(to_unsigned(43, 8)),
			1472 => std_logic_vector(to_unsigned(61, 8)),
			1473 => std_logic_vector(to_unsigned(157, 8)),
			1474 => std_logic_vector(to_unsigned(143, 8)),
			1475 => std_logic_vector(to_unsigned(145, 8)),
			1476 => std_logic_vector(to_unsigned(12, 8)),
			1477 => std_logic_vector(to_unsigned(75, 8)),
			1478 => std_logic_vector(to_unsigned(180, 8)),
			1479 => std_logic_vector(to_unsigned(237, 8)),
			1480 => std_logic_vector(to_unsigned(19, 8)),
			1481 => std_logic_vector(to_unsigned(155, 8)),
			1482 => std_logic_vector(to_unsigned(141, 8)),
			1483 => std_logic_vector(to_unsigned(238, 8)),
			1484 => std_logic_vector(to_unsigned(47, 8)),
			1485 => std_logic_vector(to_unsigned(53, 8)),
			1486 => std_logic_vector(to_unsigned(135, 8)),
			1487 => std_logic_vector(to_unsigned(218, 8)),
			1488 => std_logic_vector(to_unsigned(62, 8)),
			1489 => std_logic_vector(to_unsigned(220, 8)),
			1490 => std_logic_vector(to_unsigned(226, 8)),
			1491 => std_logic_vector(to_unsigned(170, 8)),
			1492 => std_logic_vector(to_unsigned(211, 8)),
			1493 => std_logic_vector(to_unsigned(83, 8)),
			1494 => std_logic_vector(to_unsigned(107, 8)),
			1495 => std_logic_vector(to_unsigned(220, 8)),
			1496 => std_logic_vector(to_unsigned(52, 8)),
			1497 => std_logic_vector(to_unsigned(28, 8)),
			1498 => std_logic_vector(to_unsigned(88, 8)),
			1499 => std_logic_vector(to_unsigned(251, 8)),
			1500 => std_logic_vector(to_unsigned(210, 8)),
			1501 => std_logic_vector(to_unsigned(180, 8)),
			1502 => std_logic_vector(to_unsigned(122, 8)),
			1503 => std_logic_vector(to_unsigned(181, 8)),
			1504 => std_logic_vector(to_unsigned(238, 8)),
			1505 => std_logic_vector(to_unsigned(108, 8)),
			1506 => std_logic_vector(to_unsigned(13, 8)),
			1507 => std_logic_vector(to_unsigned(41, 8)),
			1508 => std_logic_vector(to_unsigned(221, 8)),
			1509 => std_logic_vector(to_unsigned(21, 8)),
			1510 => std_logic_vector(to_unsigned(50, 8)),
			1511 => std_logic_vector(to_unsigned(109, 8)),
			1512 => std_logic_vector(to_unsigned(183, 8)),
			1513 => std_logic_vector(to_unsigned(100, 8)),
			1514 => std_logic_vector(to_unsigned(7, 8)),
			1515 => std_logic_vector(to_unsigned(209, 8)),
			1516 => std_logic_vector(to_unsigned(61, 8)),
			1517 => std_logic_vector(to_unsigned(180, 8)),
			1518 => std_logic_vector(to_unsigned(40, 8)),
			1519 => std_logic_vector(to_unsigned(31, 8)),
			1520 => std_logic_vector(to_unsigned(209, 8)),
			1521 => std_logic_vector(to_unsigned(16, 8)),
			1522 => std_logic_vector(to_unsigned(193, 8)),
			1523 => std_logic_vector(to_unsigned(241, 8)),
			1524 => std_logic_vector(to_unsigned(125, 8)),
			1525 => std_logic_vector(to_unsigned(14, 8)),
			1526 => std_logic_vector(to_unsigned(251, 8)),
			1527 => std_logic_vector(to_unsigned(20, 8)),
			1528 => std_logic_vector(to_unsigned(122, 8)),
			1529 => std_logic_vector(to_unsigned(31, 8)),
			1530 => std_logic_vector(to_unsigned(34, 8)),
			1531 => std_logic_vector(to_unsigned(61, 8)),
			1532 => std_logic_vector(to_unsigned(247, 8)),
			1533 => std_logic_vector(to_unsigned(2, 8)),
			1534 => std_logic_vector(to_unsigned(183, 8)),
			1535 => std_logic_vector(to_unsigned(167, 8)),
			1536 => std_logic_vector(to_unsigned(129, 8)),
			1537 => std_logic_vector(to_unsigned(180, 8)),
			1538 => std_logic_vector(to_unsigned(135, 8)),
			1539 => std_logic_vector(to_unsigned(103, 8)),
			1540 => std_logic_vector(to_unsigned(59, 8)),
			1541 => std_logic_vector(to_unsigned(171, 8)),
			1542 => std_logic_vector(to_unsigned(96, 8)),
			1543 => std_logic_vector(to_unsigned(113, 8)),
			1544 => std_logic_vector(to_unsigned(124, 8)),
			1545 => std_logic_vector(to_unsigned(73, 8)),
			1546 => std_logic_vector(to_unsigned(163, 8)),
			1547 => std_logic_vector(to_unsigned(10, 8)),
			1548 => std_logic_vector(to_unsigned(192, 8)),
			1549 => std_logic_vector(to_unsigned(88, 8)),
			1550 => std_logic_vector(to_unsigned(2, 8)),
			1551 => std_logic_vector(to_unsigned(75, 8)),
			1552 => std_logic_vector(to_unsigned(102, 8)),
			1553 => std_logic_vector(to_unsigned(12, 8)),
			1554 => std_logic_vector(to_unsigned(206, 8)),
			1555 => std_logic_vector(to_unsigned(73, 8)),
			1556 => std_logic_vector(to_unsigned(18, 8)),
			1557 => std_logic_vector(to_unsigned(122, 8)),
			1558 => std_logic_vector(to_unsigned(140, 8)),
			1559 => std_logic_vector(to_unsigned(201, 8)),
			1560 => std_logic_vector(to_unsigned(59, 8)),
			1561 => std_logic_vector(to_unsigned(76, 8)),
			1562 => std_logic_vector(to_unsigned(66, 8)),
			1563 => std_logic_vector(to_unsigned(175, 8)),
			1564 => std_logic_vector(to_unsigned(209, 8)),
			1565 => std_logic_vector(to_unsigned(152, 8)),
			1566 => std_logic_vector(to_unsigned(44, 8)),
			1567 => std_logic_vector(to_unsigned(197, 8)),
			1568 => std_logic_vector(to_unsigned(24, 8)),
			1569 => std_logic_vector(to_unsigned(134, 8)),
			1570 => std_logic_vector(to_unsigned(118, 8)),
			1571 => std_logic_vector(to_unsigned(120, 8)),
			1572 => std_logic_vector(to_unsigned(52, 8)),
			1573 => std_logic_vector(to_unsigned(52, 8)),
			1574 => std_logic_vector(to_unsigned(122, 8)),
			1575 => std_logic_vector(to_unsigned(115, 8)),
			1576 => std_logic_vector(to_unsigned(194, 8)),
			1577 => std_logic_vector(to_unsigned(173, 8)),
			1578 => std_logic_vector(to_unsigned(123, 8)),
			1579 => std_logic_vector(to_unsigned(16, 8)),
			1580 => std_logic_vector(to_unsigned(218, 8)),
			1581 => std_logic_vector(to_unsigned(141, 8)),
			1582 => std_logic_vector(to_unsigned(107, 8)),
			1583 => std_logic_vector(to_unsigned(6, 8)),
			1584 => std_logic_vector(to_unsigned(138, 8)),
			1585 => std_logic_vector(to_unsigned(103, 8)),
			1586 => std_logic_vector(to_unsigned(185, 8)),
			1587 => std_logic_vector(to_unsigned(54, 8)),
			1588 => std_logic_vector(to_unsigned(51, 8)),
			1589 => std_logic_vector(to_unsigned(125, 8)),
			1590 => std_logic_vector(to_unsigned(49, 8)),
			1591 => std_logic_vector(to_unsigned(255, 8)),
			1592 => std_logic_vector(to_unsigned(114, 8)),
			1593 => std_logic_vector(to_unsigned(25, 8)),
			1594 => std_logic_vector(to_unsigned(45, 8)),
			1595 => std_logic_vector(to_unsigned(31, 8)),
			1596 => std_logic_vector(to_unsigned(49, 8)),
			1597 => std_logic_vector(to_unsigned(58, 8)),
			1598 => std_logic_vector(to_unsigned(171, 8)),
			1599 => std_logic_vector(to_unsigned(153, 8)),
			1600 => std_logic_vector(to_unsigned(47, 8)),
			1601 => std_logic_vector(to_unsigned(46, 8)),
			1602 => std_logic_vector(to_unsigned(249, 8)),
			1603 => std_logic_vector(to_unsigned(11, 8)),
			1604 => std_logic_vector(to_unsigned(218, 8)),
			1605 => std_logic_vector(to_unsigned(99, 8)),
			1606 => std_logic_vector(to_unsigned(170, 8)),
			1607 => std_logic_vector(to_unsigned(58, 8)),
			1608 => std_logic_vector(to_unsigned(110, 8)),
			1609 => std_logic_vector(to_unsigned(187, 8)),
			1610 => std_logic_vector(to_unsigned(180, 8)),
			1611 => std_logic_vector(to_unsigned(170, 8)),
			1612 => std_logic_vector(to_unsigned(228, 8)),
			1613 => std_logic_vector(to_unsigned(247, 8)),
			1614 => std_logic_vector(to_unsigned(85, 8)),
			1615 => std_logic_vector(to_unsigned(191, 8)),
			1616 => std_logic_vector(to_unsigned(84, 8)),
			1617 => std_logic_vector(to_unsigned(46, 8)),
			1618 => std_logic_vector(to_unsigned(35, 8)),
			1619 => std_logic_vector(to_unsigned(180, 8)),
			1620 => std_logic_vector(to_unsigned(84, 8)),
			1621 => std_logic_vector(to_unsigned(57, 8)),
			1622 => std_logic_vector(to_unsigned(127, 8)),
			1623 => std_logic_vector(to_unsigned(232, 8)),
			1624 => std_logic_vector(to_unsigned(183, 8)),
			1625 => std_logic_vector(to_unsigned(55, 8)),
			1626 => std_logic_vector(to_unsigned(180, 8)),
			1627 => std_logic_vector(to_unsigned(22, 8)),
			1628 => std_logic_vector(to_unsigned(125, 8)),
			1629 => std_logic_vector(to_unsigned(196, 8)),
			1630 => std_logic_vector(to_unsigned(66, 8)),
			1631 => std_logic_vector(to_unsigned(19, 8)),
			1632 => std_logic_vector(to_unsigned(117, 8)),
			1633 => std_logic_vector(to_unsigned(89, 8)),
			1634 => std_logic_vector(to_unsigned(216, 8)),
			1635 => std_logic_vector(to_unsigned(43, 8)),
			1636 => std_logic_vector(to_unsigned(196, 8)),
			1637 => std_logic_vector(to_unsigned(206, 8)),
			1638 => std_logic_vector(to_unsigned(154, 8)),
			1639 => std_logic_vector(to_unsigned(209, 8)),
			1640 => std_logic_vector(to_unsigned(79, 8)),
			1641 => std_logic_vector(to_unsigned(38, 8)),
			1642 => std_logic_vector(to_unsigned(45, 8)),
			1643 => std_logic_vector(to_unsigned(6, 8)),
			1644 => std_logic_vector(to_unsigned(51, 8)),
			1645 => std_logic_vector(to_unsigned(161, 8)),
			1646 => std_logic_vector(to_unsigned(214, 8)),
			1647 => std_logic_vector(to_unsigned(253, 8)),
			1648 => std_logic_vector(to_unsigned(57, 8)),
			1649 => std_logic_vector(to_unsigned(251, 8)),
			1650 => std_logic_vector(to_unsigned(254, 8)),
			1651 => std_logic_vector(to_unsigned(165, 8)),
			1652 => std_logic_vector(to_unsigned(145, 8)),
			1653 => std_logic_vector(to_unsigned(123, 8)),
			1654 => std_logic_vector(to_unsigned(136, 8)),
			1655 => std_logic_vector(to_unsigned(39, 8)),
			1656 => std_logic_vector(to_unsigned(251, 8)),
			1657 => std_logic_vector(to_unsigned(203, 8)),
			1658 => std_logic_vector(to_unsigned(182, 8)),
			1659 => std_logic_vector(to_unsigned(127, 8)),
			1660 => std_logic_vector(to_unsigned(224, 8)),
			1661 => std_logic_vector(to_unsigned(42, 8)),
			1662 => std_logic_vector(to_unsigned(252, 8)),
			1663 => std_logic_vector(to_unsigned(80, 8)),
			1664 => std_logic_vector(to_unsigned(136, 8)),
			1665 => std_logic_vector(to_unsigned(19, 8)),
			1666 => std_logic_vector(to_unsigned(184, 8)),
			1667 => std_logic_vector(to_unsigned(33, 8)),
			1668 => std_logic_vector(to_unsigned(24, 8)),
			1669 => std_logic_vector(to_unsigned(102, 8)),
			1670 => std_logic_vector(to_unsigned(169, 8)),
			1671 => std_logic_vector(to_unsigned(178, 8)),
			1672 => std_logic_vector(to_unsigned(176, 8)),
			1673 => std_logic_vector(to_unsigned(22, 8)),
			1674 => std_logic_vector(to_unsigned(70, 8)),
			1675 => std_logic_vector(to_unsigned(119, 8)),
			1676 => std_logic_vector(to_unsigned(152, 8)),
			1677 => std_logic_vector(to_unsigned(58, 8)),
			1678 => std_logic_vector(to_unsigned(141, 8)),
			1679 => std_logic_vector(to_unsigned(97, 8)),
			1680 => std_logic_vector(to_unsigned(102, 8)),
			1681 => std_logic_vector(to_unsigned(230, 8)),
			1682 => std_logic_vector(to_unsigned(52, 8)),
			1683 => std_logic_vector(to_unsigned(204, 8)),
			1684 => std_logic_vector(to_unsigned(120, 8)),
			1685 => std_logic_vector(to_unsigned(58, 8)),
			1686 => std_logic_vector(to_unsigned(188, 8)),
			1687 => std_logic_vector(to_unsigned(211, 8)),
			1688 => std_logic_vector(to_unsigned(59, 8)),
			1689 => std_logic_vector(to_unsigned(22, 8)),
			1690 => std_logic_vector(to_unsigned(187, 8)),
			1691 => std_logic_vector(to_unsigned(23, 8)),
			1692 => std_logic_vector(to_unsigned(218, 8)),
			1693 => std_logic_vector(to_unsigned(112, 8)),
			1694 => std_logic_vector(to_unsigned(26, 8)),
			1695 => std_logic_vector(to_unsigned(123, 8)),
			1696 => std_logic_vector(to_unsigned(82, 8)),
			1697 => std_logic_vector(to_unsigned(84, 8)),
			1698 => std_logic_vector(to_unsigned(34, 8)),
			1699 => std_logic_vector(to_unsigned(203, 8)),
			1700 => std_logic_vector(to_unsigned(19, 8)),
			1701 => std_logic_vector(to_unsigned(31, 8)),
			1702 => std_logic_vector(to_unsigned(253, 8)),
			1703 => std_logic_vector(to_unsigned(35, 8)),
			1704 => std_logic_vector(to_unsigned(223, 8)),
			1705 => std_logic_vector(to_unsigned(136, 8)),
			1706 => std_logic_vector(to_unsigned(213, 8)),
			1707 => std_logic_vector(to_unsigned(27, 8)),
			1708 => std_logic_vector(to_unsigned(158, 8)),
			1709 => std_logic_vector(to_unsigned(243, 8)),
			1710 => std_logic_vector(to_unsigned(15, 8)),
			1711 => std_logic_vector(to_unsigned(13, 8)),
			1712 => std_logic_vector(to_unsigned(247, 8)),
			1713 => std_logic_vector(to_unsigned(150, 8)),
			1714 => std_logic_vector(to_unsigned(128, 8)),
			1715 => std_logic_vector(to_unsigned(216, 8)),
			1716 => std_logic_vector(to_unsigned(1, 8)),
			1717 => std_logic_vector(to_unsigned(236, 8)),
			1718 => std_logic_vector(to_unsigned(186, 8)),
			1719 => std_logic_vector(to_unsigned(212, 8)),
			1720 => std_logic_vector(to_unsigned(172, 8)),
			1721 => std_logic_vector(to_unsigned(204, 8)),
			1722 => std_logic_vector(to_unsigned(109, 8)),
			1723 => std_logic_vector(to_unsigned(119, 8)),
			others => (others => '0'));   

signal RAM1: ram_type := (0 => std_logic_vector(to_unsigned(95, 8)),
			1 => std_logic_vector(to_unsigned(38, 8)),
			2 => std_logic_vector(to_unsigned(154, 8)),
			3 => std_logic_vector(to_unsigned(5, 8)),
			4 => std_logic_vector(to_unsigned(105, 8)),
			5 => std_logic_vector(to_unsigned(177, 8)),
			6 => std_logic_vector(to_unsigned(74, 8)),
			7 => std_logic_vector(to_unsigned(129, 8)),
			8 => std_logic_vector(to_unsigned(129, 8)),
			9 => std_logic_vector(to_unsigned(60, 8)),
			10 => std_logic_vector(to_unsigned(172, 8)),
			11 => std_logic_vector(to_unsigned(99, 8)),
			12 => std_logic_vector(to_unsigned(173, 8)),
			13 => std_logic_vector(to_unsigned(99, 8)),
			14 => std_logic_vector(to_unsigned(23, 8)),
			15 => std_logic_vector(to_unsigned(69, 8)),
			16 => std_logic_vector(to_unsigned(147, 8)),
			17 => std_logic_vector(to_unsigned(249, 8)),
			18 => std_logic_vector(to_unsigned(246, 8)),
			19 => std_logic_vector(to_unsigned(192, 8)),
			20 => std_logic_vector(to_unsigned(126, 8)),
			21 => std_logic_vector(to_unsigned(210, 8)),
			22 => std_logic_vector(to_unsigned(113, 8)),
			23 => std_logic_vector(to_unsigned(213, 8)),
			24 => std_logic_vector(to_unsigned(198, 8)),
			25 => std_logic_vector(to_unsigned(71, 8)),
			26 => std_logic_vector(to_unsigned(38, 8)),
			27 => std_logic_vector(to_unsigned(167, 8)),
			28 => std_logic_vector(to_unsigned(214, 8)),
			29 => std_logic_vector(to_unsigned(138, 8)),
			30 => std_logic_vector(to_unsigned(252, 8)),
			31 => std_logic_vector(to_unsigned(116, 8)),
			32 => std_logic_vector(to_unsigned(233, 8)),
			33 => std_logic_vector(to_unsigned(12, 8)),
			34 => std_logic_vector(to_unsigned(131, 8)),
			35 => std_logic_vector(to_unsigned(183, 8)),
			36 => std_logic_vector(to_unsigned(112, 8)),
			37 => std_logic_vector(to_unsigned(255, 8)),
			38 => std_logic_vector(to_unsigned(74, 8)),
			39 => std_logic_vector(to_unsigned(127, 8)),
			40 => std_logic_vector(to_unsigned(21, 8)),
			41 => std_logic_vector(to_unsigned(161, 8)),
			42 => std_logic_vector(to_unsigned(91, 8)),
			43 => std_logic_vector(to_unsigned(142, 8)),
			44 => std_logic_vector(to_unsigned(118, 8)),
			45 => std_logic_vector(to_unsigned(30, 8)),
			46 => std_logic_vector(to_unsigned(82, 8)),
			47 => std_logic_vector(to_unsigned(143, 8)),
			48 => std_logic_vector(to_unsigned(61, 8)),
			49 => std_logic_vector(to_unsigned(160, 8)),
			50 => std_logic_vector(to_unsigned(188, 8)),
			51 => std_logic_vector(to_unsigned(34, 8)),
			52 => std_logic_vector(to_unsigned(125, 8)),
			53 => std_logic_vector(to_unsigned(220, 8)),
			54 => std_logic_vector(to_unsigned(21, 8)),
			55 => std_logic_vector(to_unsigned(126, 8)),
			56 => std_logic_vector(to_unsigned(182, 8)),
			57 => std_logic_vector(to_unsigned(20, 8)),
			58 => std_logic_vector(to_unsigned(54, 8)),
			59 => std_logic_vector(to_unsigned(240, 8)),
			60 => std_logic_vector(to_unsigned(251, 8)),
			61 => std_logic_vector(to_unsigned(182, 8)),
			62 => std_logic_vector(to_unsigned(150, 8)),
			63 => std_logic_vector(to_unsigned(15, 8)),
			64 => std_logic_vector(to_unsigned(210, 8)),
			65 => std_logic_vector(to_unsigned(202, 8)),
			66 => std_logic_vector(to_unsigned(28, 8)),
			67 => std_logic_vector(to_unsigned(1, 8)),
			68 => std_logic_vector(to_unsigned(154, 8)),
			69 => std_logic_vector(to_unsigned(150, 8)),
			70 => std_logic_vector(to_unsigned(212, 8)),
			71 => std_logic_vector(to_unsigned(44, 8)),
			72 => std_logic_vector(to_unsigned(145, 8)),
			73 => std_logic_vector(to_unsigned(117, 8)),
			74 => std_logic_vector(to_unsigned(145, 8)),
			75 => std_logic_vector(to_unsigned(26, 8)),
			76 => std_logic_vector(to_unsigned(53, 8)),
			77 => std_logic_vector(to_unsigned(21, 8)),
			78 => std_logic_vector(to_unsigned(99, 8)),
			79 => std_logic_vector(to_unsigned(13, 8)),
			80 => std_logic_vector(to_unsigned(119, 8)),
			81 => std_logic_vector(to_unsigned(124, 8)),
			82 => std_logic_vector(to_unsigned(87, 8)),
			83 => std_logic_vector(to_unsigned(249, 8)),
			84 => std_logic_vector(to_unsigned(131, 8)),
			85 => std_logic_vector(to_unsigned(78, 8)),
			86 => std_logic_vector(to_unsigned(144, 8)),
			87 => std_logic_vector(to_unsigned(152, 8)),
			88 => std_logic_vector(to_unsigned(236, 8)),
			89 => std_logic_vector(to_unsigned(247, 8)),
			90 => std_logic_vector(to_unsigned(23, 8)),
			91 => std_logic_vector(to_unsigned(51, 8)),
			92 => std_logic_vector(to_unsigned(57, 8)),
			93 => std_logic_vector(to_unsigned(245, 8)),
			94 => std_logic_vector(to_unsigned(217, 8)),
			95 => std_logic_vector(to_unsigned(106, 8)),
			96 => std_logic_vector(to_unsigned(177, 8)),
			97 => std_logic_vector(to_unsigned(189, 8)),
			98 => std_logic_vector(to_unsigned(128, 8)),
			99 => std_logic_vector(to_unsigned(31, 8)),
			100 => std_logic_vector(to_unsigned(134, 8)),
			101 => std_logic_vector(to_unsigned(103, 8)),
			102 => std_logic_vector(to_unsigned(76, 8)),
			103 => std_logic_vector(to_unsigned(167, 8)),
			104 => std_logic_vector(to_unsigned(141, 8)),
			105 => std_logic_vector(to_unsigned(209, 8)),
			106 => std_logic_vector(to_unsigned(6, 8)),
			107 => std_logic_vector(to_unsigned(61, 8)),
			108 => std_logic_vector(to_unsigned(166, 8)),
			109 => std_logic_vector(to_unsigned(150, 8)),
			110 => std_logic_vector(to_unsigned(216, 8)),
			111 => std_logic_vector(to_unsigned(102, 8)),
			112 => std_logic_vector(to_unsigned(213, 8)),
			113 => std_logic_vector(to_unsigned(183, 8)),
			114 => std_logic_vector(to_unsigned(195, 8)),
			115 => std_logic_vector(to_unsigned(234, 8)),
			116 => std_logic_vector(to_unsigned(219, 8)),
			117 => std_logic_vector(to_unsigned(24, 8)),
			118 => std_logic_vector(to_unsigned(192, 8)),
			119 => std_logic_vector(to_unsigned(105, 8)),
			120 => std_logic_vector(to_unsigned(89, 8)),
			121 => std_logic_vector(to_unsigned(93, 8)),
			122 => std_logic_vector(to_unsigned(74, 8)),
			123 => std_logic_vector(to_unsigned(28, 8)),
			124 => std_logic_vector(to_unsigned(218, 8)),
			125 => std_logic_vector(to_unsigned(197, 8)),
			126 => std_logic_vector(to_unsigned(35, 8)),
			127 => std_logic_vector(to_unsigned(187, 8)),
			128 => std_logic_vector(to_unsigned(225, 8)),
			129 => std_logic_vector(to_unsigned(103, 8)),
			130 => std_logic_vector(to_unsigned(35, 8)),
			131 => std_logic_vector(to_unsigned(43, 8)),
			132 => std_logic_vector(to_unsigned(221, 8)),
			133 => std_logic_vector(to_unsigned(107, 8)),
			134 => std_logic_vector(to_unsigned(114, 8)),
			135 => std_logic_vector(to_unsigned(73, 8)),
			136 => std_logic_vector(to_unsigned(246, 8)),
			137 => std_logic_vector(to_unsigned(241, 8)),
			138 => std_logic_vector(to_unsigned(86, 8)),
			139 => std_logic_vector(to_unsigned(137, 8)),
			140 => std_logic_vector(to_unsigned(178, 8)),
			141 => std_logic_vector(to_unsigned(145, 8)),
			142 => std_logic_vector(to_unsigned(52, 8)),
			143 => std_logic_vector(to_unsigned(228, 8)),
			144 => std_logic_vector(to_unsigned(192, 8)),
			145 => std_logic_vector(to_unsigned(170, 8)),
			146 => std_logic_vector(to_unsigned(147, 8)),
			147 => std_logic_vector(to_unsigned(31, 8)),
			148 => std_logic_vector(to_unsigned(17, 8)),
			149 => std_logic_vector(to_unsigned(244, 8)),
			150 => std_logic_vector(to_unsigned(212, 8)),
			151 => std_logic_vector(to_unsigned(28, 8)),
			152 => std_logic_vector(to_unsigned(94, 8)),
			153 => std_logic_vector(to_unsigned(224, 8)),
			154 => std_logic_vector(to_unsigned(200, 8)),
			155 => std_logic_vector(to_unsigned(224, 8)),
			156 => std_logic_vector(to_unsigned(241, 8)),
			157 => std_logic_vector(to_unsigned(15, 8)),
			158 => std_logic_vector(to_unsigned(234, 8)),
			159 => std_logic_vector(to_unsigned(41, 8)),
			160 => std_logic_vector(to_unsigned(2, 8)),
			161 => std_logic_vector(to_unsigned(87, 8)),
			162 => std_logic_vector(to_unsigned(32, 8)),
			163 => std_logic_vector(to_unsigned(7, 8)),
			164 => std_logic_vector(to_unsigned(177, 8)),
			165 => std_logic_vector(to_unsigned(139, 8)),
			166 => std_logic_vector(to_unsigned(20, 8)),
			167 => std_logic_vector(to_unsigned(136, 8)),
			168 => std_logic_vector(to_unsigned(125, 8)),
			169 => std_logic_vector(to_unsigned(186, 8)),
			170 => std_logic_vector(to_unsigned(92, 8)),
			171 => std_logic_vector(to_unsigned(163, 8)),
			172 => std_logic_vector(to_unsigned(148, 8)),
			173 => std_logic_vector(to_unsigned(139, 8)),
			174 => std_logic_vector(to_unsigned(70, 8)),
			175 => std_logic_vector(to_unsigned(184, 8)),
			176 => std_logic_vector(to_unsigned(156, 8)),
			177 => std_logic_vector(to_unsigned(115, 8)),
			178 => std_logic_vector(to_unsigned(172, 8)),
			179 => std_logic_vector(to_unsigned(164, 8)),
			180 => std_logic_vector(to_unsigned(5, 8)),
			181 => std_logic_vector(to_unsigned(71, 8)),
			182 => std_logic_vector(to_unsigned(12, 8)),
			183 => std_logic_vector(to_unsigned(204, 8)),
			184 => std_logic_vector(to_unsigned(2, 8)),
			185 => std_logic_vector(to_unsigned(14, 8)),
			186 => std_logic_vector(to_unsigned(107, 8)),
			187 => std_logic_vector(to_unsigned(103, 8)),
			188 => std_logic_vector(to_unsigned(186, 8)),
			189 => std_logic_vector(to_unsigned(134, 8)),
			190 => std_logic_vector(to_unsigned(4, 8)),
			191 => std_logic_vector(to_unsigned(205, 8)),
			192 => std_logic_vector(to_unsigned(242, 8)),
			193 => std_logic_vector(to_unsigned(113, 8)),
			194 => std_logic_vector(to_unsigned(139, 8)),
			195 => std_logic_vector(to_unsigned(37, 8)),
			196 => std_logic_vector(to_unsigned(76, 8)),
			197 => std_logic_vector(to_unsigned(23, 8)),
			198 => std_logic_vector(to_unsigned(29, 8)),
			199 => std_logic_vector(to_unsigned(20, 8)),
			200 => std_logic_vector(to_unsigned(55, 8)),
			201 => std_logic_vector(to_unsigned(118, 8)),
			202 => std_logic_vector(to_unsigned(27, 8)),
			203 => std_logic_vector(to_unsigned(182, 8)),
			204 => std_logic_vector(to_unsigned(10, 8)),
			205 => std_logic_vector(to_unsigned(0, 8)),
			206 => std_logic_vector(to_unsigned(81, 8)),
			207 => std_logic_vector(to_unsigned(134, 8)),
			208 => std_logic_vector(to_unsigned(29, 8)),
			209 => std_logic_vector(to_unsigned(248, 8)),
			210 => std_logic_vector(to_unsigned(107, 8)),
			211 => std_logic_vector(to_unsigned(110, 8)),
			212 => std_logic_vector(to_unsigned(204, 8)),
			213 => std_logic_vector(to_unsigned(174, 8)),
			214 => std_logic_vector(to_unsigned(205, 8)),
			215 => std_logic_vector(to_unsigned(179, 8)),
			216 => std_logic_vector(to_unsigned(171, 8)),
			217 => std_logic_vector(to_unsigned(130, 8)),
			218 => std_logic_vector(to_unsigned(248, 8)),
			219 => std_logic_vector(to_unsigned(48, 8)),
			220 => std_logic_vector(to_unsigned(81, 8)),
			221 => std_logic_vector(to_unsigned(198, 8)),
			222 => std_logic_vector(to_unsigned(218, 8)),
			223 => std_logic_vector(to_unsigned(206, 8)),
			224 => std_logic_vector(to_unsigned(12, 8)),
			225 => std_logic_vector(to_unsigned(136, 8)),
			226 => std_logic_vector(to_unsigned(193, 8)),
			227 => std_logic_vector(to_unsigned(82, 8)),
			228 => std_logic_vector(to_unsigned(156, 8)),
			229 => std_logic_vector(to_unsigned(10, 8)),
			230 => std_logic_vector(to_unsigned(143, 8)),
			231 => std_logic_vector(to_unsigned(228, 8)),
			232 => std_logic_vector(to_unsigned(30, 8)),
			233 => std_logic_vector(to_unsigned(191, 8)),
			234 => std_logic_vector(to_unsigned(28, 8)),
			235 => std_logic_vector(to_unsigned(116, 8)),
			236 => std_logic_vector(to_unsigned(237, 8)),
			237 => std_logic_vector(to_unsigned(16, 8)),
			238 => std_logic_vector(to_unsigned(209, 8)),
			239 => std_logic_vector(to_unsigned(209, 8)),
			240 => std_logic_vector(to_unsigned(41, 8)),
			241 => std_logic_vector(to_unsigned(106, 8)),
			242 => std_logic_vector(to_unsigned(107, 8)),
			243 => std_logic_vector(to_unsigned(145, 8)),
			244 => std_logic_vector(to_unsigned(190, 8)),
			245 => std_logic_vector(to_unsigned(173, 8)),
			246 => std_logic_vector(to_unsigned(82, 8)),
			247 => std_logic_vector(to_unsigned(33, 8)),
			248 => std_logic_vector(to_unsigned(251, 8)),
			249 => std_logic_vector(to_unsigned(69, 8)),
			250 => std_logic_vector(to_unsigned(28, 8)),
			251 => std_logic_vector(to_unsigned(75, 8)),
			252 => std_logic_vector(to_unsigned(245, 8)),
			253 => std_logic_vector(to_unsigned(151, 8)),
			254 => std_logic_vector(to_unsigned(207, 8)),
			255 => std_logic_vector(to_unsigned(75, 8)),
			256 => std_logic_vector(to_unsigned(28, 8)),
			257 => std_logic_vector(to_unsigned(238, 8)),
			258 => std_logic_vector(to_unsigned(69, 8)),
			259 => std_logic_vector(to_unsigned(118, 8)),
			260 => std_logic_vector(to_unsigned(8, 8)),
			261 => std_logic_vector(to_unsigned(12, 8)),
			262 => std_logic_vector(to_unsigned(102, 8)),
			263 => std_logic_vector(to_unsigned(89, 8)),
			264 => std_logic_vector(to_unsigned(110, 8)),
			265 => std_logic_vector(to_unsigned(44, 8)),
			266 => std_logic_vector(to_unsigned(134, 8)),
			267 => std_logic_vector(to_unsigned(254, 8)),
			268 => std_logic_vector(to_unsigned(241, 8)),
			269 => std_logic_vector(to_unsigned(165, 8)),
			270 => std_logic_vector(to_unsigned(14, 8)),
			271 => std_logic_vector(to_unsigned(21, 8)),
			272 => std_logic_vector(to_unsigned(105, 8)),
			273 => std_logic_vector(to_unsigned(156, 8)),
			274 => std_logic_vector(to_unsigned(2, 8)),
			275 => std_logic_vector(to_unsigned(57, 8)),
			276 => std_logic_vector(to_unsigned(137, 8)),
			277 => std_logic_vector(to_unsigned(101, 8)),
			278 => std_logic_vector(to_unsigned(119, 8)),
			279 => std_logic_vector(to_unsigned(151, 8)),
			280 => std_logic_vector(to_unsigned(50, 8)),
			281 => std_logic_vector(to_unsigned(35, 8)),
			282 => std_logic_vector(to_unsigned(144, 8)),
			283 => std_logic_vector(to_unsigned(8, 8)),
			284 => std_logic_vector(to_unsigned(105, 8)),
			285 => std_logic_vector(to_unsigned(208, 8)),
			286 => std_logic_vector(to_unsigned(116, 8)),
			287 => std_logic_vector(to_unsigned(153, 8)),
			288 => std_logic_vector(to_unsigned(8, 8)),
			289 => std_logic_vector(to_unsigned(109, 8)),
			290 => std_logic_vector(to_unsigned(47, 8)),
			291 => std_logic_vector(to_unsigned(13, 8)),
			292 => std_logic_vector(to_unsigned(149, 8)),
			293 => std_logic_vector(to_unsigned(127, 8)),
			294 => std_logic_vector(to_unsigned(222, 8)),
			295 => std_logic_vector(to_unsigned(185, 8)),
			296 => std_logic_vector(to_unsigned(70, 8)),
			297 => std_logic_vector(to_unsigned(207, 8)),
			298 => std_logic_vector(to_unsigned(179, 8)),
			299 => std_logic_vector(to_unsigned(6, 8)),
			300 => std_logic_vector(to_unsigned(52, 8)),
			301 => std_logic_vector(to_unsigned(79, 8)),
			302 => std_logic_vector(to_unsigned(233, 8)),
			303 => std_logic_vector(to_unsigned(180, 8)),
			304 => std_logic_vector(to_unsigned(224, 8)),
			305 => std_logic_vector(to_unsigned(44, 8)),
			306 => std_logic_vector(to_unsigned(222, 8)),
			307 => std_logic_vector(to_unsigned(130, 8)),
			308 => std_logic_vector(to_unsigned(154, 8)),
			309 => std_logic_vector(to_unsigned(9, 8)),
			310 => std_logic_vector(to_unsigned(158, 8)),
			311 => std_logic_vector(to_unsigned(147, 8)),
			312 => std_logic_vector(to_unsigned(135, 8)),
			313 => std_logic_vector(to_unsigned(170, 8)),
			314 => std_logic_vector(to_unsigned(65, 8)),
			315 => std_logic_vector(to_unsigned(104, 8)),
			316 => std_logic_vector(to_unsigned(128, 8)),
			317 => std_logic_vector(to_unsigned(45, 8)),
			318 => std_logic_vector(to_unsigned(235, 8)),
			319 => std_logic_vector(to_unsigned(126, 8)),
			320 => std_logic_vector(to_unsigned(173, 8)),
			321 => std_logic_vector(to_unsigned(253, 8)),
			322 => std_logic_vector(to_unsigned(46, 8)),
			323 => std_logic_vector(to_unsigned(28, 8)),
			324 => std_logic_vector(to_unsigned(152, 8)),
			325 => std_logic_vector(to_unsigned(126, 8)),
			326 => std_logic_vector(to_unsigned(175, 8)),
			327 => std_logic_vector(to_unsigned(233, 8)),
			328 => std_logic_vector(to_unsigned(145, 8)),
			329 => std_logic_vector(to_unsigned(95, 8)),
			330 => std_logic_vector(to_unsigned(176, 8)),
			331 => std_logic_vector(to_unsigned(91, 8)),
			332 => std_logic_vector(to_unsigned(155, 8)),
			333 => std_logic_vector(to_unsigned(207, 8)),
			334 => std_logic_vector(to_unsigned(116, 8)),
			335 => std_logic_vector(to_unsigned(60, 8)),
			336 => std_logic_vector(to_unsigned(128, 8)),
			337 => std_logic_vector(to_unsigned(209, 8)),
			338 => std_logic_vector(to_unsigned(98, 8)),
			339 => std_logic_vector(to_unsigned(128, 8)),
			340 => std_logic_vector(to_unsigned(192, 8)),
			341 => std_logic_vector(to_unsigned(209, 8)),
			342 => std_logic_vector(to_unsigned(220, 8)),
			343 => std_logic_vector(to_unsigned(254, 8)),
			344 => std_logic_vector(to_unsigned(166, 8)),
			345 => std_logic_vector(to_unsigned(165, 8)),
			346 => std_logic_vector(to_unsigned(53, 8)),
			347 => std_logic_vector(to_unsigned(93, 8)),
			348 => std_logic_vector(to_unsigned(189, 8)),
			349 => std_logic_vector(to_unsigned(4, 8)),
			350 => std_logic_vector(to_unsigned(103, 8)),
			351 => std_logic_vector(to_unsigned(181, 8)),
			352 => std_logic_vector(to_unsigned(243, 8)),
			353 => std_logic_vector(to_unsigned(136, 8)),
			354 => std_logic_vector(to_unsigned(192, 8)),
			355 => std_logic_vector(to_unsigned(135, 8)),
			356 => std_logic_vector(to_unsigned(69, 8)),
			357 => std_logic_vector(to_unsigned(84, 8)),
			358 => std_logic_vector(to_unsigned(18, 8)),
			359 => std_logic_vector(to_unsigned(99, 8)),
			360 => std_logic_vector(to_unsigned(217, 8)),
			361 => std_logic_vector(to_unsigned(99, 8)),
			362 => std_logic_vector(to_unsigned(107, 8)),
			363 => std_logic_vector(to_unsigned(172, 8)),
			364 => std_logic_vector(to_unsigned(163, 8)),
			365 => std_logic_vector(to_unsigned(100, 8)),
			366 => std_logic_vector(to_unsigned(101, 8)),
			367 => std_logic_vector(to_unsigned(246, 8)),
			368 => std_logic_vector(to_unsigned(190, 8)),
			369 => std_logic_vector(to_unsigned(122, 8)),
			370 => std_logic_vector(to_unsigned(96, 8)),
			371 => std_logic_vector(to_unsigned(89, 8)),
			372 => std_logic_vector(to_unsigned(29, 8)),
			373 => std_logic_vector(to_unsigned(181, 8)),
			374 => std_logic_vector(to_unsigned(251, 8)),
			375 => std_logic_vector(to_unsigned(206, 8)),
			376 => std_logic_vector(to_unsigned(155, 8)),
			377 => std_logic_vector(to_unsigned(205, 8)),
			378 => std_logic_vector(to_unsigned(198, 8)),
			379 => std_logic_vector(to_unsigned(131, 8)),
			380 => std_logic_vector(to_unsigned(9, 8)),
			381 => std_logic_vector(to_unsigned(241, 8)),
			382 => std_logic_vector(to_unsigned(161, 8)),
			383 => std_logic_vector(to_unsigned(122, 8)),
			384 => std_logic_vector(to_unsigned(100, 8)),
			385 => std_logic_vector(to_unsigned(184, 8)),
			386 => std_logic_vector(to_unsigned(167, 8)),
			387 => std_logic_vector(to_unsigned(36, 8)),
			388 => std_logic_vector(to_unsigned(230, 8)),
			389 => std_logic_vector(to_unsigned(160, 8)),
			390 => std_logic_vector(to_unsigned(88, 8)),
			391 => std_logic_vector(to_unsigned(35, 8)),
			392 => std_logic_vector(to_unsigned(10, 8)),
			393 => std_logic_vector(to_unsigned(122, 8)),
			394 => std_logic_vector(to_unsigned(66, 8)),
			395 => std_logic_vector(to_unsigned(155, 8)),
			396 => std_logic_vector(to_unsigned(213, 8)),
			397 => std_logic_vector(to_unsigned(6, 8)),
			398 => std_logic_vector(to_unsigned(228, 8)),
			399 => std_logic_vector(to_unsigned(12, 8)),
			400 => std_logic_vector(to_unsigned(29, 8)),
			401 => std_logic_vector(to_unsigned(225, 8)),
			402 => std_logic_vector(to_unsigned(120, 8)),
			403 => std_logic_vector(to_unsigned(155, 8)),
			404 => std_logic_vector(to_unsigned(46, 8)),
			405 => std_logic_vector(to_unsigned(43, 8)),
			406 => std_logic_vector(to_unsigned(9, 8)),
			407 => std_logic_vector(to_unsigned(34, 8)),
			408 => std_logic_vector(to_unsigned(108, 8)),
			409 => std_logic_vector(to_unsigned(132, 8)),
			410 => std_logic_vector(to_unsigned(140, 8)),
			411 => std_logic_vector(to_unsigned(61, 8)),
			412 => std_logic_vector(to_unsigned(139, 8)),
			413 => std_logic_vector(to_unsigned(222, 8)),
			414 => std_logic_vector(to_unsigned(171, 8)),
			415 => std_logic_vector(to_unsigned(82, 8)),
			416 => std_logic_vector(to_unsigned(122, 8)),
			417 => std_logic_vector(to_unsigned(42, 8)),
			418 => std_logic_vector(to_unsigned(17, 8)),
			419 => std_logic_vector(to_unsigned(189, 8)),
			420 => std_logic_vector(to_unsigned(19, 8)),
			421 => std_logic_vector(to_unsigned(128, 8)),
			422 => std_logic_vector(to_unsigned(70, 8)),
			423 => std_logic_vector(to_unsigned(248, 8)),
			424 => std_logic_vector(to_unsigned(110, 8)),
			425 => std_logic_vector(to_unsigned(107, 8)),
			426 => std_logic_vector(to_unsigned(183, 8)),
			427 => std_logic_vector(to_unsigned(108, 8)),
			428 => std_logic_vector(to_unsigned(49, 8)),
			429 => std_logic_vector(to_unsigned(22, 8)),
			430 => std_logic_vector(to_unsigned(41, 8)),
			431 => std_logic_vector(to_unsigned(131, 8)),
			432 => std_logic_vector(to_unsigned(183, 8)),
			433 => std_logic_vector(to_unsigned(9, 8)),
			434 => std_logic_vector(to_unsigned(33, 8)),
			435 => std_logic_vector(to_unsigned(152, 8)),
			436 => std_logic_vector(to_unsigned(253, 8)),
			437 => std_logic_vector(to_unsigned(68, 8)),
			438 => std_logic_vector(to_unsigned(210, 8)),
			439 => std_logic_vector(to_unsigned(201, 8)),
			440 => std_logic_vector(to_unsigned(86, 8)),
			441 => std_logic_vector(to_unsigned(77, 8)),
			442 => std_logic_vector(to_unsigned(148, 8)),
			443 => std_logic_vector(to_unsigned(247, 8)),
			444 => std_logic_vector(to_unsigned(100, 8)),
			445 => std_logic_vector(to_unsigned(26, 8)),
			446 => std_logic_vector(to_unsigned(228, 8)),
			447 => std_logic_vector(to_unsigned(47, 8)),
			448 => std_logic_vector(to_unsigned(80, 8)),
			449 => std_logic_vector(to_unsigned(219, 8)),
			450 => std_logic_vector(to_unsigned(126, 8)),
			451 => std_logic_vector(to_unsigned(85, 8)),
			452 => std_logic_vector(to_unsigned(150, 8)),
			453 => std_logic_vector(to_unsigned(57, 8)),
			454 => std_logic_vector(to_unsigned(62, 8)),
			455 => std_logic_vector(to_unsigned(53, 8)),
			456 => std_logic_vector(to_unsigned(81, 8)),
			457 => std_logic_vector(to_unsigned(254, 8)),
			458 => std_logic_vector(to_unsigned(238, 8)),
			459 => std_logic_vector(to_unsigned(192, 8)),
			460 => std_logic_vector(to_unsigned(39, 8)),
			461 => std_logic_vector(to_unsigned(57, 8)),
			462 => std_logic_vector(to_unsigned(71, 8)),
			463 => std_logic_vector(to_unsigned(111, 8)),
			464 => std_logic_vector(to_unsigned(120, 8)),
			465 => std_logic_vector(to_unsigned(205, 8)),
			466 => std_logic_vector(to_unsigned(180, 8)),
			467 => std_logic_vector(to_unsigned(247, 8)),
			468 => std_logic_vector(to_unsigned(132, 8)),
			469 => std_logic_vector(to_unsigned(33, 8)),
			470 => std_logic_vector(to_unsigned(76, 8)),
			471 => std_logic_vector(to_unsigned(231, 8)),
			472 => std_logic_vector(to_unsigned(210, 8)),
			473 => std_logic_vector(to_unsigned(110, 8)),
			474 => std_logic_vector(to_unsigned(63, 8)),
			475 => std_logic_vector(to_unsigned(16, 8)),
			476 => std_logic_vector(to_unsigned(121, 8)),
			477 => std_logic_vector(to_unsigned(154, 8)),
			478 => std_logic_vector(to_unsigned(107, 8)),
			479 => std_logic_vector(to_unsigned(126, 8)),
			480 => std_logic_vector(to_unsigned(139, 8)),
			481 => std_logic_vector(to_unsigned(103, 8)),
			482 => std_logic_vector(to_unsigned(246, 8)),
			483 => std_logic_vector(to_unsigned(29, 8)),
			484 => std_logic_vector(to_unsigned(162, 8)),
			485 => std_logic_vector(to_unsigned(0, 8)),
			486 => std_logic_vector(to_unsigned(24, 8)),
			487 => std_logic_vector(to_unsigned(107, 8)),
			488 => std_logic_vector(to_unsigned(98, 8)),
			489 => std_logic_vector(to_unsigned(218, 8)),
			490 => std_logic_vector(to_unsigned(40, 8)),
			491 => std_logic_vector(to_unsigned(243, 8)),
			492 => std_logic_vector(to_unsigned(98, 8)),
			493 => std_logic_vector(to_unsigned(240, 8)),
			494 => std_logic_vector(to_unsigned(49, 8)),
			495 => std_logic_vector(to_unsigned(191, 8)),
			496 => std_logic_vector(to_unsigned(133, 8)),
			497 => std_logic_vector(to_unsigned(114, 8)),
			498 => std_logic_vector(to_unsigned(59, 8)),
			499 => std_logic_vector(to_unsigned(193, 8)),
			500 => std_logic_vector(to_unsigned(50, 8)),
			501 => std_logic_vector(to_unsigned(147, 8)),
			502 => std_logic_vector(to_unsigned(221, 8)),
			503 => std_logic_vector(to_unsigned(110, 8)),
			504 => std_logic_vector(to_unsigned(185, 8)),
			505 => std_logic_vector(to_unsigned(217, 8)),
			506 => std_logic_vector(to_unsigned(154, 8)),
			507 => std_logic_vector(to_unsigned(227, 8)),
			508 => std_logic_vector(to_unsigned(82, 8)),
			509 => std_logic_vector(to_unsigned(127, 8)),
			510 => std_logic_vector(to_unsigned(83, 8)),
			511 => std_logic_vector(to_unsigned(122, 8)),
			512 => std_logic_vector(to_unsigned(173, 8)),
			513 => std_logic_vector(to_unsigned(35, 8)),
			514 => std_logic_vector(to_unsigned(197, 8)),
			515 => std_logic_vector(to_unsigned(92, 8)),
			516 => std_logic_vector(to_unsigned(147, 8)),
			517 => std_logic_vector(to_unsigned(71, 8)),
			518 => std_logic_vector(to_unsigned(235, 8)),
			519 => std_logic_vector(to_unsigned(88, 8)),
			520 => std_logic_vector(to_unsigned(88, 8)),
			521 => std_logic_vector(to_unsigned(80, 8)),
			522 => std_logic_vector(to_unsigned(66, 8)),
			523 => std_logic_vector(to_unsigned(62, 8)),
			524 => std_logic_vector(to_unsigned(70, 8)),
			525 => std_logic_vector(to_unsigned(165, 8)),
			526 => std_logic_vector(to_unsigned(137, 8)),
			527 => std_logic_vector(to_unsigned(13, 8)),
			528 => std_logic_vector(to_unsigned(143, 8)),
			529 => std_logic_vector(to_unsigned(196, 8)),
			530 => std_logic_vector(to_unsigned(98, 8)),
			531 => std_logic_vector(to_unsigned(117, 8)),
			532 => std_logic_vector(to_unsigned(108, 8)),
			533 => std_logic_vector(to_unsigned(144, 8)),
			534 => std_logic_vector(to_unsigned(85, 8)),
			535 => std_logic_vector(to_unsigned(224, 8)),
			536 => std_logic_vector(to_unsigned(190, 8)),
			537 => std_logic_vector(to_unsigned(181, 8)),
			538 => std_logic_vector(to_unsigned(252, 8)),
			539 => std_logic_vector(to_unsigned(135, 8)),
			540 => std_logic_vector(to_unsigned(96, 8)),
			541 => std_logic_vector(to_unsigned(95, 8)),
			542 => std_logic_vector(to_unsigned(17, 8)),
			543 => std_logic_vector(to_unsigned(22, 8)),
			544 => std_logic_vector(to_unsigned(26, 8)),
			545 => std_logic_vector(to_unsigned(181, 8)),
			546 => std_logic_vector(to_unsigned(133, 8)),
			547 => std_logic_vector(to_unsigned(255, 8)),
			548 => std_logic_vector(to_unsigned(134, 8)),
			549 => std_logic_vector(to_unsigned(175, 8)),
			550 => std_logic_vector(to_unsigned(91, 8)),
			551 => std_logic_vector(to_unsigned(22, 8)),
			552 => std_logic_vector(to_unsigned(58, 8)),
			553 => std_logic_vector(to_unsigned(193, 8)),
			554 => std_logic_vector(to_unsigned(200, 8)),
			555 => std_logic_vector(to_unsigned(252, 8)),
			556 => std_logic_vector(to_unsigned(115, 8)),
			557 => std_logic_vector(to_unsigned(54, 8)),
			558 => std_logic_vector(to_unsigned(227, 8)),
			559 => std_logic_vector(to_unsigned(232, 8)),
			560 => std_logic_vector(to_unsigned(163, 8)),
			561 => std_logic_vector(to_unsigned(216, 8)),
			562 => std_logic_vector(to_unsigned(60, 8)),
			563 => std_logic_vector(to_unsigned(165, 8)),
			564 => std_logic_vector(to_unsigned(54, 8)),
			565 => std_logic_vector(to_unsigned(250, 8)),
			566 => std_logic_vector(to_unsigned(201, 8)),
			567 => std_logic_vector(to_unsigned(27, 8)),
			568 => std_logic_vector(to_unsigned(139, 8)),
			569 => std_logic_vector(to_unsigned(62, 8)),
			570 => std_logic_vector(to_unsigned(166, 8)),
			571 => std_logic_vector(to_unsigned(121, 8)),
			572 => std_logic_vector(to_unsigned(48, 8)),
			573 => std_logic_vector(to_unsigned(167, 8)),
			574 => std_logic_vector(to_unsigned(92, 8)),
			575 => std_logic_vector(to_unsigned(89, 8)),
			576 => std_logic_vector(to_unsigned(254, 8)),
			577 => std_logic_vector(to_unsigned(19, 8)),
			578 => std_logic_vector(to_unsigned(234, 8)),
			579 => std_logic_vector(to_unsigned(180, 8)),
			580 => std_logic_vector(to_unsigned(147, 8)),
			581 => std_logic_vector(to_unsigned(221, 8)),
			582 => std_logic_vector(to_unsigned(18, 8)),
			583 => std_logic_vector(to_unsigned(22, 8)),
			584 => std_logic_vector(to_unsigned(197, 8)),
			585 => std_logic_vector(to_unsigned(29, 8)),
			586 => std_logic_vector(to_unsigned(73, 8)),
			587 => std_logic_vector(to_unsigned(95, 8)),
			588 => std_logic_vector(to_unsigned(37, 8)),
			589 => std_logic_vector(to_unsigned(234, 8)),
			590 => std_logic_vector(to_unsigned(73, 8)),
			591 => std_logic_vector(to_unsigned(81, 8)),
			592 => std_logic_vector(to_unsigned(79, 8)),
			593 => std_logic_vector(to_unsigned(178, 8)),
			594 => std_logic_vector(to_unsigned(2, 8)),
			595 => std_logic_vector(to_unsigned(93, 8)),
			596 => std_logic_vector(to_unsigned(135, 8)),
			597 => std_logic_vector(to_unsigned(41, 8)),
			598 => std_logic_vector(to_unsigned(118, 8)),
			599 => std_logic_vector(to_unsigned(81, 8)),
			600 => std_logic_vector(to_unsigned(55, 8)),
			601 => std_logic_vector(to_unsigned(248, 8)),
			602 => std_logic_vector(to_unsigned(55, 8)),
			603 => std_logic_vector(to_unsigned(166, 8)),
			604 => std_logic_vector(to_unsigned(143, 8)),
			605 => std_logic_vector(to_unsigned(234, 8)),
			606 => std_logic_vector(to_unsigned(103, 8)),
			607 => std_logic_vector(to_unsigned(112, 8)),
			608 => std_logic_vector(to_unsigned(183, 8)),
			609 => std_logic_vector(to_unsigned(143, 8)),
			610 => std_logic_vector(to_unsigned(238, 8)),
			611 => std_logic_vector(to_unsigned(125, 8)),
			612 => std_logic_vector(to_unsigned(234, 8)),
			613 => std_logic_vector(to_unsigned(137, 8)),
			614 => std_logic_vector(to_unsigned(21, 8)),
			615 => std_logic_vector(to_unsigned(95, 8)),
			616 => std_logic_vector(to_unsigned(184, 8)),
			617 => std_logic_vector(to_unsigned(51, 8)),
			618 => std_logic_vector(to_unsigned(75, 8)),
			619 => std_logic_vector(to_unsigned(152, 8)),
			620 => std_logic_vector(to_unsigned(78, 8)),
			621 => std_logic_vector(to_unsigned(176, 8)),
			622 => std_logic_vector(to_unsigned(78, 8)),
			623 => std_logic_vector(to_unsigned(199, 8)),
			624 => std_logic_vector(to_unsigned(218, 8)),
			625 => std_logic_vector(to_unsigned(75, 8)),
			626 => std_logic_vector(to_unsigned(140, 8)),
			627 => std_logic_vector(to_unsigned(120, 8)),
			628 => std_logic_vector(to_unsigned(210, 8)),
			629 => std_logic_vector(to_unsigned(214, 8)),
			630 => std_logic_vector(to_unsigned(110, 8)),
			631 => std_logic_vector(to_unsigned(139, 8)),
			632 => std_logic_vector(to_unsigned(128, 8)),
			633 => std_logic_vector(to_unsigned(64, 8)),
			634 => std_logic_vector(to_unsigned(147, 8)),
			635 => std_logic_vector(to_unsigned(228, 8)),
			636 => std_logic_vector(to_unsigned(172, 8)),
			637 => std_logic_vector(to_unsigned(188, 8)),
			638 => std_logic_vector(to_unsigned(5, 8)),
			639 => std_logic_vector(to_unsigned(180, 8)),
			640 => std_logic_vector(to_unsigned(216, 8)),
			641 => std_logic_vector(to_unsigned(23, 8)),
			642 => std_logic_vector(to_unsigned(127, 8)),
			643 => std_logic_vector(to_unsigned(116, 8)),
			644 => std_logic_vector(to_unsigned(178, 8)),
			645 => std_logic_vector(to_unsigned(225, 8)),
			646 => std_logic_vector(to_unsigned(211, 8)),
			647 => std_logic_vector(to_unsigned(203, 8)),
			648 => std_logic_vector(to_unsigned(72, 8)),
			649 => std_logic_vector(to_unsigned(59, 8)),
			650 => std_logic_vector(to_unsigned(222, 8)),
			651 => std_logic_vector(to_unsigned(103, 8)),
			652 => std_logic_vector(to_unsigned(166, 8)),
			653 => std_logic_vector(to_unsigned(190, 8)),
			654 => std_logic_vector(to_unsigned(19, 8)),
			655 => std_logic_vector(to_unsigned(66, 8)),
			656 => std_logic_vector(to_unsigned(142, 8)),
			657 => std_logic_vector(to_unsigned(181, 8)),
			658 => std_logic_vector(to_unsigned(48, 8)),
			659 => std_logic_vector(to_unsigned(175, 8)),
			660 => std_logic_vector(to_unsigned(33, 8)),
			661 => std_logic_vector(to_unsigned(164, 8)),
			662 => std_logic_vector(to_unsigned(99, 8)),
			663 => std_logic_vector(to_unsigned(144, 8)),
			664 => std_logic_vector(to_unsigned(61, 8)),
			665 => std_logic_vector(to_unsigned(71, 8)),
			666 => std_logic_vector(to_unsigned(195, 8)),
			667 => std_logic_vector(to_unsigned(78, 8)),
			668 => std_logic_vector(to_unsigned(82, 8)),
			669 => std_logic_vector(to_unsigned(56, 8)),
			670 => std_logic_vector(to_unsigned(80, 8)),
			671 => std_logic_vector(to_unsigned(13, 8)),
			672 => std_logic_vector(to_unsigned(82, 8)),
			673 => std_logic_vector(to_unsigned(46, 8)),
			674 => std_logic_vector(to_unsigned(150, 8)),
			675 => std_logic_vector(to_unsigned(94, 8)),
			676 => std_logic_vector(to_unsigned(131, 8)),
			677 => std_logic_vector(to_unsigned(252, 8)),
			678 => std_logic_vector(to_unsigned(77, 8)),
			679 => std_logic_vector(to_unsigned(18, 8)),
			680 => std_logic_vector(to_unsigned(97, 8)),
			681 => std_logic_vector(to_unsigned(128, 8)),
			682 => std_logic_vector(to_unsigned(141, 8)),
			683 => std_logic_vector(to_unsigned(94, 8)),
			684 => std_logic_vector(to_unsigned(81, 8)),
			685 => std_logic_vector(to_unsigned(12, 8)),
			686 => std_logic_vector(to_unsigned(144, 8)),
			687 => std_logic_vector(to_unsigned(104, 8)),
			688 => std_logic_vector(to_unsigned(127, 8)),
			689 => std_logic_vector(to_unsigned(65, 8)),
			690 => std_logic_vector(to_unsigned(58, 8)),
			691 => std_logic_vector(to_unsigned(89, 8)),
			692 => std_logic_vector(to_unsigned(166, 8)),
			693 => std_logic_vector(to_unsigned(106, 8)),
			694 => std_logic_vector(to_unsigned(119, 8)),
			695 => std_logic_vector(to_unsigned(95, 8)),
			696 => std_logic_vector(to_unsigned(195, 8)),
			697 => std_logic_vector(to_unsigned(71, 8)),
			698 => std_logic_vector(to_unsigned(106, 8)),
			699 => std_logic_vector(to_unsigned(113, 8)),
			700 => std_logic_vector(to_unsigned(204, 8)),
			701 => std_logic_vector(to_unsigned(62, 8)),
			702 => std_logic_vector(to_unsigned(239, 8)),
			703 => std_logic_vector(to_unsigned(167, 8)),
			704 => std_logic_vector(to_unsigned(250, 8)),
			705 => std_logic_vector(to_unsigned(11, 8)),
			706 => std_logic_vector(to_unsigned(234, 8)),
			707 => std_logic_vector(to_unsigned(221, 8)),
			708 => std_logic_vector(to_unsigned(86, 8)),
			709 => std_logic_vector(to_unsigned(149, 8)),
			710 => std_logic_vector(to_unsigned(253, 8)),
			711 => std_logic_vector(to_unsigned(239, 8)),
			712 => std_logic_vector(to_unsigned(32, 8)),
			713 => std_logic_vector(to_unsigned(20, 8)),
			714 => std_logic_vector(to_unsigned(26, 8)),
			715 => std_logic_vector(to_unsigned(137, 8)),
			716 => std_logic_vector(to_unsigned(238, 8)),
			717 => std_logic_vector(to_unsigned(37, 8)),
			718 => std_logic_vector(to_unsigned(54, 8)),
			719 => std_logic_vector(to_unsigned(145, 8)),
			720 => std_logic_vector(to_unsigned(55, 8)),
			721 => std_logic_vector(to_unsigned(48, 8)),
			722 => std_logic_vector(to_unsigned(82, 8)),
			723 => std_logic_vector(to_unsigned(120, 8)),
			724 => std_logic_vector(to_unsigned(187, 8)),
			725 => std_logic_vector(to_unsigned(85, 8)),
			726 => std_logic_vector(to_unsigned(197, 8)),
			727 => std_logic_vector(to_unsigned(167, 8)),
			728 => std_logic_vector(to_unsigned(124, 8)),
			729 => std_logic_vector(to_unsigned(231, 8)),
			730 => std_logic_vector(to_unsigned(181, 8)),
			731 => std_logic_vector(to_unsigned(15, 8)),
			732 => std_logic_vector(to_unsigned(250, 8)),
			733 => std_logic_vector(to_unsigned(218, 8)),
			734 => std_logic_vector(to_unsigned(247, 8)),
			735 => std_logic_vector(to_unsigned(128, 8)),
			736 => std_logic_vector(to_unsigned(231, 8)),
			737 => std_logic_vector(to_unsigned(190, 8)),
			738 => std_logic_vector(to_unsigned(213, 8)),
			739 => std_logic_vector(to_unsigned(247, 8)),
			740 => std_logic_vector(to_unsigned(107, 8)),
			741 => std_logic_vector(to_unsigned(56, 8)),
			742 => std_logic_vector(to_unsigned(250, 8)),
			743 => std_logic_vector(to_unsigned(100, 8)),
			744 => std_logic_vector(to_unsigned(83, 8)),
			745 => std_logic_vector(to_unsigned(47, 8)),
			746 => std_logic_vector(to_unsigned(166, 8)),
			747 => std_logic_vector(to_unsigned(16, 8)),
			748 => std_logic_vector(to_unsigned(56, 8)),
			749 => std_logic_vector(to_unsigned(42, 8)),
			750 => std_logic_vector(to_unsigned(223, 8)),
			751 => std_logic_vector(to_unsigned(192, 8)),
			752 => std_logic_vector(to_unsigned(229, 8)),
			753 => std_logic_vector(to_unsigned(193, 8)),
			754 => std_logic_vector(to_unsigned(116, 8)),
			755 => std_logic_vector(to_unsigned(42, 8)),
			756 => std_logic_vector(to_unsigned(104, 8)),
			757 => std_logic_vector(to_unsigned(131, 8)),
			758 => std_logic_vector(to_unsigned(54, 8)),
			759 => std_logic_vector(to_unsigned(148, 8)),
			760 => std_logic_vector(to_unsigned(138, 8)),
			761 => std_logic_vector(to_unsigned(222, 8)),
			762 => std_logic_vector(to_unsigned(3, 8)),
			763 => std_logic_vector(to_unsigned(184, 8)),
			764 => std_logic_vector(to_unsigned(230, 8)),
			765 => std_logic_vector(to_unsigned(33, 8)),
			766 => std_logic_vector(to_unsigned(231, 8)),
			767 => std_logic_vector(to_unsigned(169, 8)),
			768 => std_logic_vector(to_unsigned(52, 8)),
			769 => std_logic_vector(to_unsigned(133, 8)),
			770 => std_logic_vector(to_unsigned(117, 8)),
			771 => std_logic_vector(to_unsigned(183, 8)),
			772 => std_logic_vector(to_unsigned(176, 8)),
			773 => std_logic_vector(to_unsigned(192, 8)),
			774 => std_logic_vector(to_unsigned(225, 8)),
			775 => std_logic_vector(to_unsigned(245, 8)),
			776 => std_logic_vector(to_unsigned(151, 8)),
			777 => std_logic_vector(to_unsigned(201, 8)),
			778 => std_logic_vector(to_unsigned(142, 8)),
			779 => std_logic_vector(to_unsigned(23, 8)),
			780 => std_logic_vector(to_unsigned(135, 8)),
			781 => std_logic_vector(to_unsigned(241, 8)),
			782 => std_logic_vector(to_unsigned(212, 8)),
			783 => std_logic_vector(to_unsigned(54, 8)),
			784 => std_logic_vector(to_unsigned(92, 8)),
			785 => std_logic_vector(to_unsigned(106, 8)),
			786 => std_logic_vector(to_unsigned(98, 8)),
			787 => std_logic_vector(to_unsigned(97, 8)),
			788 => std_logic_vector(to_unsigned(226, 8)),
			789 => std_logic_vector(to_unsigned(245, 8)),
			790 => std_logic_vector(to_unsigned(87, 8)),
			791 => std_logic_vector(to_unsigned(59, 8)),
			792 => std_logic_vector(to_unsigned(70, 8)),
			793 => std_logic_vector(to_unsigned(229, 8)),
			794 => std_logic_vector(to_unsigned(7, 8)),
			795 => std_logic_vector(to_unsigned(127, 8)),
			796 => std_logic_vector(to_unsigned(179, 8)),
			797 => std_logic_vector(to_unsigned(100, 8)),
			798 => std_logic_vector(to_unsigned(170, 8)),
			799 => std_logic_vector(to_unsigned(68, 8)),
			800 => std_logic_vector(to_unsigned(44, 8)),
			801 => std_logic_vector(to_unsigned(18, 8)),
			802 => std_logic_vector(to_unsigned(95, 8)),
			803 => std_logic_vector(to_unsigned(114, 8)),
			804 => std_logic_vector(to_unsigned(151, 8)),
			805 => std_logic_vector(to_unsigned(211, 8)),
			806 => std_logic_vector(to_unsigned(51, 8)),
			807 => std_logic_vector(to_unsigned(149, 8)),
			808 => std_logic_vector(to_unsigned(175, 8)),
			809 => std_logic_vector(to_unsigned(126, 8)),
			810 => std_logic_vector(to_unsigned(201, 8)),
			811 => std_logic_vector(to_unsigned(129, 8)),
			812 => std_logic_vector(to_unsigned(7, 8)),
			813 => std_logic_vector(to_unsigned(8, 8)),
			814 => std_logic_vector(to_unsigned(254, 8)),
			815 => std_logic_vector(to_unsigned(142, 8)),
			816 => std_logic_vector(to_unsigned(146, 8)),
			817 => std_logic_vector(to_unsigned(211, 8)),
			818 => std_logic_vector(to_unsigned(141, 8)),
			819 => std_logic_vector(to_unsigned(41, 8)),
			820 => std_logic_vector(to_unsigned(71, 8)),
			821 => std_logic_vector(to_unsigned(0, 8)),
			822 => std_logic_vector(to_unsigned(137, 8)),
			823 => std_logic_vector(to_unsigned(232, 8)),
			824 => std_logic_vector(to_unsigned(40, 8)),
			825 => std_logic_vector(to_unsigned(219, 8)),
			826 => std_logic_vector(to_unsigned(129, 8)),
			827 => std_logic_vector(to_unsigned(155, 8)),
			828 => std_logic_vector(to_unsigned(113, 8)),
			829 => std_logic_vector(to_unsigned(84, 8)),
			830 => std_logic_vector(to_unsigned(93, 8)),
			831 => std_logic_vector(to_unsigned(162, 8)),
			832 => std_logic_vector(to_unsigned(188, 8)),
			833 => std_logic_vector(to_unsigned(96, 8)),
			834 => std_logic_vector(to_unsigned(173, 8)),
			835 => std_logic_vector(to_unsigned(21, 8)),
			836 => std_logic_vector(to_unsigned(49, 8)),
			837 => std_logic_vector(to_unsigned(251, 8)),
			838 => std_logic_vector(to_unsigned(255, 8)),
			839 => std_logic_vector(to_unsigned(129, 8)),
			840 => std_logic_vector(to_unsigned(51, 8)),
			841 => std_logic_vector(to_unsigned(55, 8)),
			842 => std_logic_vector(to_unsigned(124, 8)),
			843 => std_logic_vector(to_unsigned(45, 8)),
			844 => std_logic_vector(to_unsigned(202, 8)),
			845 => std_logic_vector(to_unsigned(188, 8)),
			846 => std_logic_vector(to_unsigned(91, 8)),
			847 => std_logic_vector(to_unsigned(174, 8)),
			848 => std_logic_vector(to_unsigned(168, 8)),
			849 => std_logic_vector(to_unsigned(134, 8)),
			850 => std_logic_vector(to_unsigned(160, 8)),
			851 => std_logic_vector(to_unsigned(145, 8)),
			852 => std_logic_vector(to_unsigned(84, 8)),
			853 => std_logic_vector(to_unsigned(197, 8)),
			854 => std_logic_vector(to_unsigned(16, 8)),
			855 => std_logic_vector(to_unsigned(209, 8)),
			856 => std_logic_vector(to_unsigned(129, 8)),
			857 => std_logic_vector(to_unsigned(224, 8)),
			858 => std_logic_vector(to_unsigned(173, 8)),
			859 => std_logic_vector(to_unsigned(178, 8)),
			860 => std_logic_vector(to_unsigned(98, 8)),
			861 => std_logic_vector(to_unsigned(124, 8)),
			862 => std_logic_vector(to_unsigned(252, 8)),
			863 => std_logic_vector(to_unsigned(213, 8)),
			864 => std_logic_vector(to_unsigned(27, 8)),
			865 => std_logic_vector(to_unsigned(247, 8)),
			866 => std_logic_vector(to_unsigned(103, 8)),
			867 => std_logic_vector(to_unsigned(2, 8)),
			868 => std_logic_vector(to_unsigned(121, 8)),
			869 => std_logic_vector(to_unsigned(181, 8)),
			870 => std_logic_vector(to_unsigned(84, 8)),
			871 => std_logic_vector(to_unsigned(41, 8)),
			872 => std_logic_vector(to_unsigned(146, 8)),
			873 => std_logic_vector(to_unsigned(189, 8)),
			874 => std_logic_vector(to_unsigned(12, 8)),
			875 => std_logic_vector(to_unsigned(190, 8)),
			876 => std_logic_vector(to_unsigned(71, 8)),
			877 => std_logic_vector(to_unsigned(29, 8)),
			878 => std_logic_vector(to_unsigned(205, 8)),
			879 => std_logic_vector(to_unsigned(151, 8)),
			880 => std_logic_vector(to_unsigned(239, 8)),
			881 => std_logic_vector(to_unsigned(121, 8)),
			882 => std_logic_vector(to_unsigned(222, 8)),
			883 => std_logic_vector(to_unsigned(192, 8)),
			884 => std_logic_vector(to_unsigned(231, 8)),
			885 => std_logic_vector(to_unsigned(146, 8)),
			886 => std_logic_vector(to_unsigned(46, 8)),
			887 => std_logic_vector(to_unsigned(178, 8)),
			888 => std_logic_vector(to_unsigned(35, 8)),
			889 => std_logic_vector(to_unsigned(10, 8)),
			890 => std_logic_vector(to_unsigned(154, 8)),
			891 => std_logic_vector(to_unsigned(218, 8)),
			892 => std_logic_vector(to_unsigned(239, 8)),
			893 => std_logic_vector(to_unsigned(44, 8)),
			894 => std_logic_vector(to_unsigned(67, 8)),
			895 => std_logic_vector(to_unsigned(223, 8)),
			896 => std_logic_vector(to_unsigned(196, 8)),
			897 => std_logic_vector(to_unsigned(206, 8)),
			898 => std_logic_vector(to_unsigned(166, 8)),
			899 => std_logic_vector(to_unsigned(149, 8)),
			900 => std_logic_vector(to_unsigned(33, 8)),
			901 => std_logic_vector(to_unsigned(218, 8)),
			902 => std_logic_vector(to_unsigned(123, 8)),
			903 => std_logic_vector(to_unsigned(65, 8)),
			904 => std_logic_vector(to_unsigned(52, 8)),
			905 => std_logic_vector(to_unsigned(65, 8)),
			906 => std_logic_vector(to_unsigned(85, 8)),
			907 => std_logic_vector(to_unsigned(133, 8)),
			908 => std_logic_vector(to_unsigned(26, 8)),
			909 => std_logic_vector(to_unsigned(75, 8)),
			910 => std_logic_vector(to_unsigned(110, 8)),
			911 => std_logic_vector(to_unsigned(115, 8)),
			912 => std_logic_vector(to_unsigned(16, 8)),
			913 => std_logic_vector(to_unsigned(56, 8)),
			914 => std_logic_vector(to_unsigned(56, 8)),
			915 => std_logic_vector(to_unsigned(59, 8)),
			916 => std_logic_vector(to_unsigned(116, 8)),
			917 => std_logic_vector(to_unsigned(64, 8)),
			918 => std_logic_vector(to_unsigned(209, 8)),
			919 => std_logic_vector(to_unsigned(178, 8)),
			920 => std_logic_vector(to_unsigned(162, 8)),
			921 => std_logic_vector(to_unsigned(81, 8)),
			922 => std_logic_vector(to_unsigned(87, 8)),
			923 => std_logic_vector(to_unsigned(40, 8)),
			924 => std_logic_vector(to_unsigned(205, 8)),
			925 => std_logic_vector(to_unsigned(172, 8)),
			926 => std_logic_vector(to_unsigned(7, 8)),
			927 => std_logic_vector(to_unsigned(160, 8)),
			928 => std_logic_vector(to_unsigned(168, 8)),
			929 => std_logic_vector(to_unsigned(55, 8)),
			930 => std_logic_vector(to_unsigned(29, 8)),
			931 => std_logic_vector(to_unsigned(70, 8)),
			932 => std_logic_vector(to_unsigned(198, 8)),
			933 => std_logic_vector(to_unsigned(88, 8)),
			934 => std_logic_vector(to_unsigned(105, 8)),
			935 => std_logic_vector(to_unsigned(208, 8)),
			936 => std_logic_vector(to_unsigned(0, 8)),
			937 => std_logic_vector(to_unsigned(190, 8)),
			938 => std_logic_vector(to_unsigned(206, 8)),
			939 => std_logic_vector(to_unsigned(138, 8)),
			940 => std_logic_vector(to_unsigned(2, 8)),
			941 => std_logic_vector(to_unsigned(199, 8)),
			942 => std_logic_vector(to_unsigned(19, 8)),
			943 => std_logic_vector(to_unsigned(10, 8)),
			944 => std_logic_vector(to_unsigned(120, 8)),
			945 => std_logic_vector(to_unsigned(199, 8)),
			946 => std_logic_vector(to_unsigned(7, 8)),
			947 => std_logic_vector(to_unsigned(142, 8)),
			948 => std_logic_vector(to_unsigned(248, 8)),
			949 => std_logic_vector(to_unsigned(180, 8)),
			950 => std_logic_vector(to_unsigned(14, 8)),
			951 => std_logic_vector(to_unsigned(12, 8)),
			952 => std_logic_vector(to_unsigned(178, 8)),
			953 => std_logic_vector(to_unsigned(135, 8)),
			954 => std_logic_vector(to_unsigned(25, 8)),
			955 => std_logic_vector(to_unsigned(166, 8)),
			956 => std_logic_vector(to_unsigned(97, 8)),
			957 => std_logic_vector(to_unsigned(139, 8)),
			958 => std_logic_vector(to_unsigned(207, 8)),
			959 => std_logic_vector(to_unsigned(97, 8)),
			960 => std_logic_vector(to_unsigned(63, 8)),
			961 => std_logic_vector(to_unsigned(218, 8)),
			962 => std_logic_vector(to_unsigned(16, 8)),
			963 => std_logic_vector(to_unsigned(149, 8)),
			964 => std_logic_vector(to_unsigned(250, 8)),
			965 => std_logic_vector(to_unsigned(111, 8)),
			966 => std_logic_vector(to_unsigned(78, 8)),
			967 => std_logic_vector(to_unsigned(235, 8)),
			968 => std_logic_vector(to_unsigned(255, 8)),
			969 => std_logic_vector(to_unsigned(115, 8)),
			970 => std_logic_vector(to_unsigned(23, 8)),
			971 => std_logic_vector(to_unsigned(208, 8)),
			972 => std_logic_vector(to_unsigned(21, 8)),
			973 => std_logic_vector(to_unsigned(217, 8)),
			974 => std_logic_vector(to_unsigned(237, 8)),
			975 => std_logic_vector(to_unsigned(217, 8)),
			976 => std_logic_vector(to_unsigned(155, 8)),
			977 => std_logic_vector(to_unsigned(126, 8)),
			978 => std_logic_vector(to_unsigned(100, 8)),
			979 => std_logic_vector(to_unsigned(240, 8)),
			980 => std_logic_vector(to_unsigned(70, 8)),
			981 => std_logic_vector(to_unsigned(185, 8)),
			982 => std_logic_vector(to_unsigned(11, 8)),
			983 => std_logic_vector(to_unsigned(244, 8)),
			984 => std_logic_vector(to_unsigned(253, 8)),
			985 => std_logic_vector(to_unsigned(251, 8)),
			986 => std_logic_vector(to_unsigned(240, 8)),
			987 => std_logic_vector(to_unsigned(168, 8)),
			988 => std_logic_vector(to_unsigned(193, 8)),
			989 => std_logic_vector(to_unsigned(114, 8)),
			990 => std_logic_vector(to_unsigned(229, 8)),
			991 => std_logic_vector(to_unsigned(223, 8)),
			992 => std_logic_vector(to_unsigned(168, 8)),
			993 => std_logic_vector(to_unsigned(185, 8)),
			994 => std_logic_vector(to_unsigned(221, 8)),
			995 => std_logic_vector(to_unsigned(204, 8)),
			996 => std_logic_vector(to_unsigned(42, 8)),
			997 => std_logic_vector(to_unsigned(71, 8)),
			998 => std_logic_vector(to_unsigned(227, 8)),
			999 => std_logic_vector(to_unsigned(85, 8)),
			1000 => std_logic_vector(to_unsigned(45, 8)),
			1001 => std_logic_vector(to_unsigned(158, 8)),
			1002 => std_logic_vector(to_unsigned(110, 8)),
			1003 => std_logic_vector(to_unsigned(163, 8)),
			1004 => std_logic_vector(to_unsigned(152, 8)),
			1005 => std_logic_vector(to_unsigned(80, 8)),
			1006 => std_logic_vector(to_unsigned(67, 8)),
			1007 => std_logic_vector(to_unsigned(114, 8)),
			1008 => std_logic_vector(to_unsigned(174, 8)),
			1009 => std_logic_vector(to_unsigned(138, 8)),
			1010 => std_logic_vector(to_unsigned(165, 8)),
			1011 => std_logic_vector(to_unsigned(228, 8)),
			1012 => std_logic_vector(to_unsigned(169, 8)),
			1013 => std_logic_vector(to_unsigned(17, 8)),
			1014 => std_logic_vector(to_unsigned(186, 8)),
			1015 => std_logic_vector(to_unsigned(38, 8)),
			1016 => std_logic_vector(to_unsigned(62, 8)),
			1017 => std_logic_vector(to_unsigned(67, 8)),
			1018 => std_logic_vector(to_unsigned(66, 8)),
			1019 => std_logic_vector(to_unsigned(176, 8)),
			1020 => std_logic_vector(to_unsigned(83, 8)),
			1021 => std_logic_vector(to_unsigned(252, 8)),
			1022 => std_logic_vector(to_unsigned(168, 8)),
			1023 => std_logic_vector(to_unsigned(251, 8)),
			1024 => std_logic_vector(to_unsigned(15, 8)),
			1025 => std_logic_vector(to_unsigned(208, 8)),
			1026 => std_logic_vector(to_unsigned(29, 8)),
			1027 => std_logic_vector(to_unsigned(117, 8)),
			1028 => std_logic_vector(to_unsigned(74, 8)),
			1029 => std_logic_vector(to_unsigned(25, 8)),
			1030 => std_logic_vector(to_unsigned(195, 8)),
			1031 => std_logic_vector(to_unsigned(168, 8)),
			1032 => std_logic_vector(to_unsigned(49, 8)),
			1033 => std_logic_vector(to_unsigned(193, 8)),
			1034 => std_logic_vector(to_unsigned(214, 8)),
			1035 => std_logic_vector(to_unsigned(194, 8)),
			1036 => std_logic_vector(to_unsigned(29, 8)),
			1037 => std_logic_vector(to_unsigned(211, 8)),
			1038 => std_logic_vector(to_unsigned(130, 8)),
			1039 => std_logic_vector(to_unsigned(227, 8)),
			1040 => std_logic_vector(to_unsigned(0, 8)),
			1041 => std_logic_vector(to_unsigned(139, 8)),
			1042 => std_logic_vector(to_unsigned(13, 8)),
			1043 => std_logic_vector(to_unsigned(180, 8)),
			1044 => std_logic_vector(to_unsigned(19, 8)),
			1045 => std_logic_vector(to_unsigned(193, 8)),
			1046 => std_logic_vector(to_unsigned(58, 8)),
			1047 => std_logic_vector(to_unsigned(35, 8)),
			1048 => std_logic_vector(to_unsigned(239, 8)),
			1049 => std_logic_vector(to_unsigned(133, 8)),
			1050 => std_logic_vector(to_unsigned(202, 8)),
			1051 => std_logic_vector(to_unsigned(253, 8)),
			1052 => std_logic_vector(to_unsigned(221, 8)),
			1053 => std_logic_vector(to_unsigned(0, 8)),
			1054 => std_logic_vector(to_unsigned(16, 8)),
			1055 => std_logic_vector(to_unsigned(52, 8)),
			1056 => std_logic_vector(to_unsigned(216, 8)),
			1057 => std_logic_vector(to_unsigned(21, 8)),
			1058 => std_logic_vector(to_unsigned(7, 8)),
			1059 => std_logic_vector(to_unsigned(147, 8)),
			1060 => std_logic_vector(to_unsigned(108, 8)),
			1061 => std_logic_vector(to_unsigned(241, 8)),
			1062 => std_logic_vector(to_unsigned(185, 8)),
			1063 => std_logic_vector(to_unsigned(229, 8)),
			1064 => std_logic_vector(to_unsigned(83, 8)),
			1065 => std_logic_vector(to_unsigned(218, 8)),
			1066 => std_logic_vector(to_unsigned(199, 8)),
			1067 => std_logic_vector(to_unsigned(52, 8)),
			1068 => std_logic_vector(to_unsigned(50, 8)),
			1069 => std_logic_vector(to_unsigned(85, 8)),
			1070 => std_logic_vector(to_unsigned(61, 8)),
			1071 => std_logic_vector(to_unsigned(187, 8)),
			1072 => std_logic_vector(to_unsigned(118, 8)),
			1073 => std_logic_vector(to_unsigned(232, 8)),
			1074 => std_logic_vector(to_unsigned(234, 8)),
			1075 => std_logic_vector(to_unsigned(242, 8)),
			1076 => std_logic_vector(to_unsigned(251, 8)),
			1077 => std_logic_vector(to_unsigned(51, 8)),
			1078 => std_logic_vector(to_unsigned(5, 8)),
			1079 => std_logic_vector(to_unsigned(69, 8)),
			1080 => std_logic_vector(to_unsigned(124, 8)),
			1081 => std_logic_vector(to_unsigned(169, 8)),
			1082 => std_logic_vector(to_unsigned(219, 8)),
			1083 => std_logic_vector(to_unsigned(110, 8)),
			1084 => std_logic_vector(to_unsigned(23, 8)),
			1085 => std_logic_vector(to_unsigned(28, 8)),
			1086 => std_logic_vector(to_unsigned(56, 8)),
			1087 => std_logic_vector(to_unsigned(25, 8)),
			1088 => std_logic_vector(to_unsigned(79, 8)),
			1089 => std_logic_vector(to_unsigned(176, 8)),
			1090 => std_logic_vector(to_unsigned(14, 8)),
			1091 => std_logic_vector(to_unsigned(91, 8)),
			1092 => std_logic_vector(to_unsigned(95, 8)),
			1093 => std_logic_vector(to_unsigned(222, 8)),
			1094 => std_logic_vector(to_unsigned(88, 8)),
			1095 => std_logic_vector(to_unsigned(168, 8)),
			1096 => std_logic_vector(to_unsigned(61, 8)),
			1097 => std_logic_vector(to_unsigned(10, 8)),
			1098 => std_logic_vector(to_unsigned(127, 8)),
			1099 => std_logic_vector(to_unsigned(96, 8)),
			1100 => std_logic_vector(to_unsigned(225, 8)),
			1101 => std_logic_vector(to_unsigned(166, 8)),
			1102 => std_logic_vector(to_unsigned(149, 8)),
			1103 => std_logic_vector(to_unsigned(167, 8)),
			1104 => std_logic_vector(to_unsigned(135, 8)),
			1105 => std_logic_vector(to_unsigned(58, 8)),
			1106 => std_logic_vector(to_unsigned(164, 8)),
			1107 => std_logic_vector(to_unsigned(6, 8)),
			1108 => std_logic_vector(to_unsigned(255, 8)),
			1109 => std_logic_vector(to_unsigned(56, 8)),
			1110 => std_logic_vector(to_unsigned(121, 8)),
			1111 => std_logic_vector(to_unsigned(119, 8)),
			1112 => std_logic_vector(to_unsigned(210, 8)),
			1113 => std_logic_vector(to_unsigned(201, 8)),
			1114 => std_logic_vector(to_unsigned(115, 8)),
			1115 => std_logic_vector(to_unsigned(8, 8)),
			1116 => std_logic_vector(to_unsigned(222, 8)),
			1117 => std_logic_vector(to_unsigned(148, 8)),
			1118 => std_logic_vector(to_unsigned(75, 8)),
			1119 => std_logic_vector(to_unsigned(143, 8)),
			1120 => std_logic_vector(to_unsigned(219, 8)),
			1121 => std_logic_vector(to_unsigned(94, 8)),
			1122 => std_logic_vector(to_unsigned(175, 8)),
			1123 => std_logic_vector(to_unsigned(1, 8)),
			1124 => std_logic_vector(to_unsigned(242, 8)),
			1125 => std_logic_vector(to_unsigned(112, 8)),
			1126 => std_logic_vector(to_unsigned(121, 8)),
			1127 => std_logic_vector(to_unsigned(185, 8)),
			1128 => std_logic_vector(to_unsigned(101, 8)),
			1129 => std_logic_vector(to_unsigned(34, 8)),
			1130 => std_logic_vector(to_unsigned(28, 8)),
			1131 => std_logic_vector(to_unsigned(221, 8)),
			1132 => std_logic_vector(to_unsigned(198, 8)),
			1133 => std_logic_vector(to_unsigned(52, 8)),
			1134 => std_logic_vector(to_unsigned(255, 8)),
			1135 => std_logic_vector(to_unsigned(72, 8)),
			1136 => std_logic_vector(to_unsigned(164, 8)),
			1137 => std_logic_vector(to_unsigned(56, 8)),
			1138 => std_logic_vector(to_unsigned(44, 8)),
			1139 => std_logic_vector(to_unsigned(170, 8)),
			1140 => std_logic_vector(to_unsigned(203, 8)),
			1141 => std_logic_vector(to_unsigned(88, 8)),
			1142 => std_logic_vector(to_unsigned(10, 8)),
			1143 => std_logic_vector(to_unsigned(195, 8)),
			1144 => std_logic_vector(to_unsigned(186, 8)),
			1145 => std_logic_vector(to_unsigned(155, 8)),
			1146 => std_logic_vector(to_unsigned(93, 8)),
			1147 => std_logic_vector(to_unsigned(26, 8)),
			1148 => std_logic_vector(to_unsigned(174, 8)),
			1149 => std_logic_vector(to_unsigned(195, 8)),
			1150 => std_logic_vector(to_unsigned(26, 8)),
			1151 => std_logic_vector(to_unsigned(157, 8)),
			1152 => std_logic_vector(to_unsigned(129, 8)),
			1153 => std_logic_vector(to_unsigned(153, 8)),
			1154 => std_logic_vector(to_unsigned(45, 8)),
			1155 => std_logic_vector(to_unsigned(85, 8)),
			1156 => std_logic_vector(to_unsigned(202, 8)),
			1157 => std_logic_vector(to_unsigned(119, 8)),
			1158 => std_logic_vector(to_unsigned(140, 8)),
			1159 => std_logic_vector(to_unsigned(103, 8)),
			1160 => std_logic_vector(to_unsigned(98, 8)),
			1161 => std_logic_vector(to_unsigned(185, 8)),
			1162 => std_logic_vector(to_unsigned(234, 8)),
			1163 => std_logic_vector(to_unsigned(157, 8)),
			1164 => std_logic_vector(to_unsigned(194, 8)),
			1165 => std_logic_vector(to_unsigned(15, 8)),
			1166 => std_logic_vector(to_unsigned(140, 8)),
			1167 => std_logic_vector(to_unsigned(205, 8)),
			1168 => std_logic_vector(to_unsigned(1, 8)),
			1169 => std_logic_vector(to_unsigned(132, 8)),
			1170 => std_logic_vector(to_unsigned(97, 8)),
			1171 => std_logic_vector(to_unsigned(64, 8)),
			1172 => std_logic_vector(to_unsigned(204, 8)),
			1173 => std_logic_vector(to_unsigned(194, 8)),
			1174 => std_logic_vector(to_unsigned(86, 8)),
			1175 => std_logic_vector(to_unsigned(232, 8)),
			1176 => std_logic_vector(to_unsigned(160, 8)),
			1177 => std_logic_vector(to_unsigned(241, 8)),
			1178 => std_logic_vector(to_unsigned(185, 8)),
			1179 => std_logic_vector(to_unsigned(164, 8)),
			1180 => std_logic_vector(to_unsigned(114, 8)),
			1181 => std_logic_vector(to_unsigned(24, 8)),
			1182 => std_logic_vector(to_unsigned(96, 8)),
			1183 => std_logic_vector(to_unsigned(76, 8)),
			1184 => std_logic_vector(to_unsigned(236, 8)),
			1185 => std_logic_vector(to_unsigned(50, 8)),
			1186 => std_logic_vector(to_unsigned(121, 8)),
			1187 => std_logic_vector(to_unsigned(208, 8)),
			1188 => std_logic_vector(to_unsigned(22, 8)),
			1189 => std_logic_vector(to_unsigned(249, 8)),
			1190 => std_logic_vector(to_unsigned(251, 8)),
			1191 => std_logic_vector(to_unsigned(24, 8)),
			1192 => std_logic_vector(to_unsigned(12, 8)),
			1193 => std_logic_vector(to_unsigned(181, 8)),
			1194 => std_logic_vector(to_unsigned(72, 8)),
			1195 => std_logic_vector(to_unsigned(11, 8)),
			1196 => std_logic_vector(to_unsigned(71, 8)),
			1197 => std_logic_vector(to_unsigned(151, 8)),
			1198 => std_logic_vector(to_unsigned(53, 8)),
			1199 => std_logic_vector(to_unsigned(151, 8)),
			1200 => std_logic_vector(to_unsigned(39, 8)),
			1201 => std_logic_vector(to_unsigned(73, 8)),
			1202 => std_logic_vector(to_unsigned(246, 8)),
			1203 => std_logic_vector(to_unsigned(136, 8)),
			1204 => std_logic_vector(to_unsigned(83, 8)),
			1205 => std_logic_vector(to_unsigned(150, 8)),
			1206 => std_logic_vector(to_unsigned(242, 8)),
			1207 => std_logic_vector(to_unsigned(200, 8)),
			1208 => std_logic_vector(to_unsigned(83, 8)),
			1209 => std_logic_vector(to_unsigned(157, 8)),
			1210 => std_logic_vector(to_unsigned(43, 8)),
			1211 => std_logic_vector(to_unsigned(82, 8)),
			1212 => std_logic_vector(to_unsigned(230, 8)),
			1213 => std_logic_vector(to_unsigned(107, 8)),
			1214 => std_logic_vector(to_unsigned(42, 8)),
			1215 => std_logic_vector(to_unsigned(153, 8)),
			1216 => std_logic_vector(to_unsigned(187, 8)),
			1217 => std_logic_vector(to_unsigned(183, 8)),
			1218 => std_logic_vector(to_unsigned(43, 8)),
			1219 => std_logic_vector(to_unsigned(65, 8)),
			1220 => std_logic_vector(to_unsigned(186, 8)),
			1221 => std_logic_vector(to_unsigned(124, 8)),
			1222 => std_logic_vector(to_unsigned(38, 8)),
			1223 => std_logic_vector(to_unsigned(80, 8)),
			1224 => std_logic_vector(to_unsigned(199, 8)),
			1225 => std_logic_vector(to_unsigned(110, 8)),
			1226 => std_logic_vector(to_unsigned(217, 8)),
			1227 => std_logic_vector(to_unsigned(174, 8)),
			1228 => std_logic_vector(to_unsigned(251, 8)),
			1229 => std_logic_vector(to_unsigned(142, 8)),
			1230 => std_logic_vector(to_unsigned(239, 8)),
			1231 => std_logic_vector(to_unsigned(211, 8)),
			1232 => std_logic_vector(to_unsigned(145, 8)),
			1233 => std_logic_vector(to_unsigned(43, 8)),
			1234 => std_logic_vector(to_unsigned(107, 8)),
			1235 => std_logic_vector(to_unsigned(210, 8)),
			1236 => std_logic_vector(to_unsigned(96, 8)),
			1237 => std_logic_vector(to_unsigned(125, 8)),
			1238 => std_logic_vector(to_unsigned(35, 8)),
			1239 => std_logic_vector(to_unsigned(223, 8)),
			1240 => std_logic_vector(to_unsigned(194, 8)),
			1241 => std_logic_vector(to_unsigned(27, 8)),
			1242 => std_logic_vector(to_unsigned(43, 8)),
			1243 => std_logic_vector(to_unsigned(184, 8)),
			1244 => std_logic_vector(to_unsigned(15, 8)),
			1245 => std_logic_vector(to_unsigned(51, 8)),
			1246 => std_logic_vector(to_unsigned(157, 8)),
			1247 => std_logic_vector(to_unsigned(187, 8)),
			1248 => std_logic_vector(to_unsigned(138, 8)),
			1249 => std_logic_vector(to_unsigned(92, 8)),
			1250 => std_logic_vector(to_unsigned(85, 8)),
			1251 => std_logic_vector(to_unsigned(64, 8)),
			1252 => std_logic_vector(to_unsigned(38, 8)),
			1253 => std_logic_vector(to_unsigned(159, 8)),
			1254 => std_logic_vector(to_unsigned(50, 8)),
			1255 => std_logic_vector(to_unsigned(27, 8)),
			1256 => std_logic_vector(to_unsigned(172, 8)),
			1257 => std_logic_vector(to_unsigned(82, 8)),
			1258 => std_logic_vector(to_unsigned(61, 8)),
			1259 => std_logic_vector(to_unsigned(115, 8)),
			1260 => std_logic_vector(to_unsigned(173, 8)),
			1261 => std_logic_vector(to_unsigned(73, 8)),
			1262 => std_logic_vector(to_unsigned(147, 8)),
			1263 => std_logic_vector(to_unsigned(245, 8)),
			1264 => std_logic_vector(to_unsigned(186, 8)),
			1265 => std_logic_vector(to_unsigned(243, 8)),
			1266 => std_logic_vector(to_unsigned(163, 8)),
			1267 => std_logic_vector(to_unsigned(124, 8)),
			1268 => std_logic_vector(to_unsigned(226, 8)),
			1269 => std_logic_vector(to_unsigned(39, 8)),
			1270 => std_logic_vector(to_unsigned(185, 8)),
			1271 => std_logic_vector(to_unsigned(182, 8)),
			1272 => std_logic_vector(to_unsigned(247, 8)),
			1273 => std_logic_vector(to_unsigned(212, 8)),
			1274 => std_logic_vector(to_unsigned(39, 8)),
			1275 => std_logic_vector(to_unsigned(217, 8)),
			1276 => std_logic_vector(to_unsigned(79, 8)),
			1277 => std_logic_vector(to_unsigned(244, 8)),
			1278 => std_logic_vector(to_unsigned(107, 8)),
			1279 => std_logic_vector(to_unsigned(137, 8)),
			1280 => std_logic_vector(to_unsigned(196, 8)),
			1281 => std_logic_vector(to_unsigned(254, 8)),
			1282 => std_logic_vector(to_unsigned(103, 8)),
			1283 => std_logic_vector(to_unsigned(67, 8)),
			1284 => std_logic_vector(to_unsigned(137, 8)),
			1285 => std_logic_vector(to_unsigned(155, 8)),
			1286 => std_logic_vector(to_unsigned(128, 8)),
			1287 => std_logic_vector(to_unsigned(212, 8)),
			1288 => std_logic_vector(to_unsigned(9, 8)),
			1289 => std_logic_vector(to_unsigned(57, 8)),
			1290 => std_logic_vector(to_unsigned(237, 8)),
			1291 => std_logic_vector(to_unsigned(195, 8)),
			1292 => std_logic_vector(to_unsigned(211, 8)),
			1293 => std_logic_vector(to_unsigned(253, 8)),
			1294 => std_logic_vector(to_unsigned(3, 8)),
			1295 => std_logic_vector(to_unsigned(163, 8)),
			1296 => std_logic_vector(to_unsigned(0, 8)),
			1297 => std_logic_vector(to_unsigned(234, 8)),
			1298 => std_logic_vector(to_unsigned(210, 8)),
			1299 => std_logic_vector(to_unsigned(186, 8)),
			1300 => std_logic_vector(to_unsigned(171, 8)),
			1301 => std_logic_vector(to_unsigned(247, 8)),
			1302 => std_logic_vector(to_unsigned(116, 8)),
			1303 => std_logic_vector(to_unsigned(34, 8)),
			1304 => std_logic_vector(to_unsigned(134, 8)),
			1305 => std_logic_vector(to_unsigned(154, 8)),
			1306 => std_logic_vector(to_unsigned(109, 8)),
			1307 => std_logic_vector(to_unsigned(109, 8)),
			1308 => std_logic_vector(to_unsigned(136, 8)),
			1309 => std_logic_vector(to_unsigned(9, 8)),
			1310 => std_logic_vector(to_unsigned(215, 8)),
			1311 => std_logic_vector(to_unsigned(150, 8)),
			1312 => std_logic_vector(to_unsigned(104, 8)),
			1313 => std_logic_vector(to_unsigned(112, 8)),
			1314 => std_logic_vector(to_unsigned(7, 8)),
			1315 => std_logic_vector(to_unsigned(35, 8)),
			1316 => std_logic_vector(to_unsigned(81, 8)),
			1317 => std_logic_vector(to_unsigned(212, 8)),
			1318 => std_logic_vector(to_unsigned(192, 8)),
			1319 => std_logic_vector(to_unsigned(209, 8)),
			1320 => std_logic_vector(to_unsigned(53, 8)),
			1321 => std_logic_vector(to_unsigned(223, 8)),
			1322 => std_logic_vector(to_unsigned(37, 8)),
			1323 => std_logic_vector(to_unsigned(158, 8)),
			1324 => std_logic_vector(to_unsigned(25, 8)),
			1325 => std_logic_vector(to_unsigned(137, 8)),
			1326 => std_logic_vector(to_unsigned(193, 8)),
			1327 => std_logic_vector(to_unsigned(75, 8)),
			1328 => std_logic_vector(to_unsigned(115, 8)),
			1329 => std_logic_vector(to_unsigned(69, 8)),
			1330 => std_logic_vector(to_unsigned(234, 8)),
			1331 => std_logic_vector(to_unsigned(51, 8)),
			1332 => std_logic_vector(to_unsigned(93, 8)),
			1333 => std_logic_vector(to_unsigned(187, 8)),
			1334 => std_logic_vector(to_unsigned(80, 8)),
			1335 => std_logic_vector(to_unsigned(54, 8)),
			1336 => std_logic_vector(to_unsigned(158, 8)),
			1337 => std_logic_vector(to_unsigned(240, 8)),
			1338 => std_logic_vector(to_unsigned(88, 8)),
			1339 => std_logic_vector(to_unsigned(203, 8)),
			1340 => std_logic_vector(to_unsigned(191, 8)),
			1341 => std_logic_vector(to_unsigned(90, 8)),
			1342 => std_logic_vector(to_unsigned(73, 8)),
			1343 => std_logic_vector(to_unsigned(38, 8)),
			1344 => std_logic_vector(to_unsigned(244, 8)),
			1345 => std_logic_vector(to_unsigned(24, 8)),
			1346 => std_logic_vector(to_unsigned(64, 8)),
			1347 => std_logic_vector(to_unsigned(91, 8)),
			1348 => std_logic_vector(to_unsigned(81, 8)),
			1349 => std_logic_vector(to_unsigned(158, 8)),
			1350 => std_logic_vector(to_unsigned(144, 8)),
			1351 => std_logic_vector(to_unsigned(94, 8)),
			1352 => std_logic_vector(to_unsigned(167, 8)),
			1353 => std_logic_vector(to_unsigned(232, 8)),
			1354 => std_logic_vector(to_unsigned(17, 8)),
			1355 => std_logic_vector(to_unsigned(144, 8)),
			1356 => std_logic_vector(to_unsigned(223, 8)),
			1357 => std_logic_vector(to_unsigned(33, 8)),
			1358 => std_logic_vector(to_unsigned(127, 8)),
			1359 => std_logic_vector(to_unsigned(134, 8)),
			1360 => std_logic_vector(to_unsigned(245, 8)),
			1361 => std_logic_vector(to_unsigned(43, 8)),
			1362 => std_logic_vector(to_unsigned(0, 8)),
			1363 => std_logic_vector(to_unsigned(226, 8)),
			1364 => std_logic_vector(to_unsigned(192, 8)),
			1365 => std_logic_vector(to_unsigned(43, 8)),
			1366 => std_logic_vector(to_unsigned(213, 8)),
			1367 => std_logic_vector(to_unsigned(212, 8)),
			1368 => std_logic_vector(to_unsigned(237, 8)),
			1369 => std_logic_vector(to_unsigned(149, 8)),
			1370 => std_logic_vector(to_unsigned(149, 8)),
			1371 => std_logic_vector(to_unsigned(232, 8)),
			1372 => std_logic_vector(to_unsigned(235, 8)),
			1373 => std_logic_vector(to_unsigned(6, 8)),
			1374 => std_logic_vector(to_unsigned(5, 8)),
			1375 => std_logic_vector(to_unsigned(188, 8)),
			1376 => std_logic_vector(to_unsigned(118, 8)),
			1377 => std_logic_vector(to_unsigned(199, 8)),
			1378 => std_logic_vector(to_unsigned(64, 8)),
			1379 => std_logic_vector(to_unsigned(111, 8)),
			1380 => std_logic_vector(to_unsigned(20, 8)),
			1381 => std_logic_vector(to_unsigned(35, 8)),
			1382 => std_logic_vector(to_unsigned(35, 8)),
			1383 => std_logic_vector(to_unsigned(248, 8)),
			1384 => std_logic_vector(to_unsigned(42, 8)),
			1385 => std_logic_vector(to_unsigned(12, 8)),
			1386 => std_logic_vector(to_unsigned(179, 8)),
			1387 => std_logic_vector(to_unsigned(14, 8)),
			1388 => std_logic_vector(to_unsigned(171, 8)),
			1389 => std_logic_vector(to_unsigned(178, 8)),
			1390 => std_logic_vector(to_unsigned(176, 8)),
			1391 => std_logic_vector(to_unsigned(48, 8)),
			1392 => std_logic_vector(to_unsigned(133, 8)),
			1393 => std_logic_vector(to_unsigned(241, 8)),
			1394 => std_logic_vector(to_unsigned(26, 8)),
			1395 => std_logic_vector(to_unsigned(244, 8)),
			1396 => std_logic_vector(to_unsigned(64, 8)),
			1397 => std_logic_vector(to_unsigned(134, 8)),
			1398 => std_logic_vector(to_unsigned(52, 8)),
			1399 => std_logic_vector(to_unsigned(250, 8)),
			1400 => std_logic_vector(to_unsigned(63, 8)),
			1401 => std_logic_vector(to_unsigned(16, 8)),
			1402 => std_logic_vector(to_unsigned(168, 8)),
			1403 => std_logic_vector(to_unsigned(152, 8)),
			1404 => std_logic_vector(to_unsigned(206, 8)),
			1405 => std_logic_vector(to_unsigned(87, 8)),
			1406 => std_logic_vector(to_unsigned(166, 8)),
			1407 => std_logic_vector(to_unsigned(150, 8)),
			1408 => std_logic_vector(to_unsigned(250, 8)),
			1409 => std_logic_vector(to_unsigned(81, 8)),
			1410 => std_logic_vector(to_unsigned(146, 8)),
			1411 => std_logic_vector(to_unsigned(52, 8)),
			1412 => std_logic_vector(to_unsigned(213, 8)),
			1413 => std_logic_vector(to_unsigned(227, 8)),
			1414 => std_logic_vector(to_unsigned(147, 8)),
			1415 => std_logic_vector(to_unsigned(245, 8)),
			1416 => std_logic_vector(to_unsigned(52, 8)),
			1417 => std_logic_vector(to_unsigned(175, 8)),
			1418 => std_logic_vector(to_unsigned(183, 8)),
			1419 => std_logic_vector(to_unsigned(119, 8)),
			1420 => std_logic_vector(to_unsigned(218, 8)),
			1421 => std_logic_vector(to_unsigned(235, 8)),
			1422 => std_logic_vector(to_unsigned(210, 8)),
			1423 => std_logic_vector(to_unsigned(199, 8)),
			1424 => std_logic_vector(to_unsigned(82, 8)),
			1425 => std_logic_vector(to_unsigned(199, 8)),
			1426 => std_logic_vector(to_unsigned(72, 8)),
			1427 => std_logic_vector(to_unsigned(149, 8)),
			1428 => std_logic_vector(to_unsigned(158, 8)),
			1429 => std_logic_vector(to_unsigned(13, 8)),
			1430 => std_logic_vector(to_unsigned(186, 8)),
			1431 => std_logic_vector(to_unsigned(27, 8)),
			1432 => std_logic_vector(to_unsigned(57, 8)),
			1433 => std_logic_vector(to_unsigned(184, 8)),
			1434 => std_logic_vector(to_unsigned(66, 8)),
			1435 => std_logic_vector(to_unsigned(171, 8)),
			1436 => std_logic_vector(to_unsigned(207, 8)),
			1437 => std_logic_vector(to_unsigned(151, 8)),
			1438 => std_logic_vector(to_unsigned(7, 8)),
			1439 => std_logic_vector(to_unsigned(103, 8)),
			1440 => std_logic_vector(to_unsigned(69, 8)),
			1441 => std_logic_vector(to_unsigned(39, 8)),
			1442 => std_logic_vector(to_unsigned(13, 8)),
			1443 => std_logic_vector(to_unsigned(170, 8)),
			1444 => std_logic_vector(to_unsigned(121, 8)),
			1445 => std_logic_vector(to_unsigned(250, 8)),
			1446 => std_logic_vector(to_unsigned(166, 8)),
			1447 => std_logic_vector(to_unsigned(124, 8)),
			1448 => std_logic_vector(to_unsigned(113, 8)),
			1449 => std_logic_vector(to_unsigned(210, 8)),
			1450 => std_logic_vector(to_unsigned(105, 8)),
			1451 => std_logic_vector(to_unsigned(17, 8)),
			1452 => std_logic_vector(to_unsigned(92, 8)),
			1453 => std_logic_vector(to_unsigned(209, 8)),
			1454 => std_logic_vector(to_unsigned(214, 8)),
			1455 => std_logic_vector(to_unsigned(37, 8)),
			1456 => std_logic_vector(to_unsigned(155, 8)),
			1457 => std_logic_vector(to_unsigned(177, 8)),
			1458 => std_logic_vector(to_unsigned(101, 8)),
			1459 => std_logic_vector(to_unsigned(15, 8)),
			1460 => std_logic_vector(to_unsigned(218, 8)),
			1461 => std_logic_vector(to_unsigned(103, 8)),
			1462 => std_logic_vector(to_unsigned(240, 8)),
			1463 => std_logic_vector(to_unsigned(26, 8)),
			1464 => std_logic_vector(to_unsigned(59, 8)),
			1465 => std_logic_vector(to_unsigned(200, 8)),
			1466 => std_logic_vector(to_unsigned(82, 8)),
			1467 => std_logic_vector(to_unsigned(182, 8)),
			1468 => std_logic_vector(to_unsigned(15, 8)),
			1469 => std_logic_vector(to_unsigned(166, 8)),
			1470 => std_logic_vector(to_unsigned(43, 8)),
			1471 => std_logic_vector(to_unsigned(225, 8)),
			1472 => std_logic_vector(to_unsigned(246, 8)),
			1473 => std_logic_vector(to_unsigned(6, 8)),
			1474 => std_logic_vector(to_unsigned(198, 8)),
			1475 => std_logic_vector(to_unsigned(140, 8)),
			1476 => std_logic_vector(to_unsigned(238, 8)),
			1477 => std_logic_vector(to_unsigned(230, 8)),
			1478 => std_logic_vector(to_unsigned(242, 8)),
			1479 => std_logic_vector(to_unsigned(14, 8)),
			1480 => std_logic_vector(to_unsigned(85, 8)),
			1481 => std_logic_vector(to_unsigned(77, 8)),
			1482 => std_logic_vector(to_unsigned(229, 8)),
			1483 => std_logic_vector(to_unsigned(11, 8)),
			1484 => std_logic_vector(to_unsigned(147, 8)),
			1485 => std_logic_vector(to_unsigned(143, 8)),
			1486 => std_logic_vector(to_unsigned(148, 8)),
			1487 => std_logic_vector(to_unsigned(62, 8)),
			1488 => std_logic_vector(to_unsigned(151, 8)),
			1489 => std_logic_vector(to_unsigned(109, 8)),
			1490 => std_logic_vector(to_unsigned(85, 8)),
			1491 => std_logic_vector(to_unsigned(217, 8)),
			1492 => std_logic_vector(to_unsigned(70, 8)),
			1493 => std_logic_vector(to_unsigned(120, 8)),
			1494 => std_logic_vector(to_unsigned(59, 8)),
			1495 => std_logic_vector(to_unsigned(217, 8)),
			1496 => std_logic_vector(to_unsigned(109, 8)),
			1497 => std_logic_vector(to_unsigned(251, 8)),
			1498 => std_logic_vector(to_unsigned(225, 8)),
			1499 => std_logic_vector(to_unsigned(126, 8)),
			1500 => std_logic_vector(to_unsigned(76, 8)),
			1501 => std_logic_vector(to_unsigned(90, 8)),
			1502 => std_logic_vector(to_unsigned(201, 8)),
			1503 => std_logic_vector(to_unsigned(123, 8)),
			1504 => std_logic_vector(to_unsigned(157, 8)),
			1505 => std_logic_vector(to_unsigned(223, 8)),
			1506 => std_logic_vector(to_unsigned(209, 8)),
			1507 => std_logic_vector(to_unsigned(89, 8)),
			1508 => std_logic_vector(to_unsigned(147, 8)),
			1509 => std_logic_vector(to_unsigned(187, 8)),
			1510 => std_logic_vector(to_unsigned(56, 8)),
			1511 => std_logic_vector(to_unsigned(246, 8)),
			1512 => std_logic_vector(to_unsigned(6, 8)),
			1513 => std_logic_vector(to_unsigned(26, 8)),
			1514 => std_logic_vector(to_unsigned(134, 8)),
			1515 => std_logic_vector(to_unsigned(254, 8)),
			1516 => std_logic_vector(to_unsigned(78, 8)),
			1517 => std_logic_vector(to_unsigned(117, 8)),
			1518 => std_logic_vector(to_unsigned(210, 8)),
			1519 => std_logic_vector(to_unsigned(235, 8)),
			1520 => std_logic_vector(to_unsigned(234, 8)),
			1521 => std_logic_vector(to_unsigned(243, 8)),
			1522 => std_logic_vector(to_unsigned(173, 8)),
			1523 => std_logic_vector(to_unsigned(55, 8)),
			1524 => std_logic_vector(to_unsigned(101, 8)),
			1525 => std_logic_vector(to_unsigned(85, 8)),
			1526 => std_logic_vector(to_unsigned(121, 8)),
			1527 => std_logic_vector(to_unsigned(189, 8)),
			1528 => std_logic_vector(to_unsigned(250, 8)),
			1529 => std_logic_vector(to_unsigned(148, 8)),
			1530 => std_logic_vector(to_unsigned(124, 8)),
			1531 => std_logic_vector(to_unsigned(20, 8)),
			1532 => std_logic_vector(to_unsigned(194, 8)),
			1533 => std_logic_vector(to_unsigned(78, 8)),
			1534 => std_logic_vector(to_unsigned(9, 8)),
			1535 => std_logic_vector(to_unsigned(52, 8)),
			1536 => std_logic_vector(to_unsigned(207, 8)),
			1537 => std_logic_vector(to_unsigned(195, 8)),
			1538 => std_logic_vector(to_unsigned(162, 8)),
			1539 => std_logic_vector(to_unsigned(202, 8)),
			1540 => std_logic_vector(to_unsigned(248, 8)),
			1541 => std_logic_vector(to_unsigned(231, 8)),
			1542 => std_logic_vector(to_unsigned(236, 8)),
			1543 => std_logic_vector(to_unsigned(232, 8)),
			1544 => std_logic_vector(to_unsigned(79, 8)),
			1545 => std_logic_vector(to_unsigned(229, 8)),
			1546 => std_logic_vector(to_unsigned(210, 8)),
			1547 => std_logic_vector(to_unsigned(131, 8)),
			1548 => std_logic_vector(to_unsigned(228, 8)),
			1549 => std_logic_vector(to_unsigned(24, 8)),
			1550 => std_logic_vector(to_unsigned(116, 8)),
			1551 => std_logic_vector(to_unsigned(210, 8)),
			1552 => std_logic_vector(to_unsigned(104, 8)),
			1553 => std_logic_vector(to_unsigned(120, 8)),
			1554 => std_logic_vector(to_unsigned(86, 8)),
			1555 => std_logic_vector(to_unsigned(74, 8)),
			1556 => std_logic_vector(to_unsigned(42, 8)),
			1557 => std_logic_vector(to_unsigned(240, 8)),
			1558 => std_logic_vector(to_unsigned(130, 8)),
			1559 => std_logic_vector(to_unsigned(253, 8)),
			1560 => std_logic_vector(to_unsigned(44, 8)),
			1561 => std_logic_vector(to_unsigned(50, 8)),
			1562 => std_logic_vector(to_unsigned(238, 8)),
			1563 => std_logic_vector(to_unsigned(45, 8)),
			1564 => std_logic_vector(to_unsigned(138, 8)),
			1565 => std_logic_vector(to_unsigned(26, 8)),
			1566 => std_logic_vector(to_unsigned(43, 8)),
			1567 => std_logic_vector(to_unsigned(77, 8)),
			1568 => std_logic_vector(to_unsigned(71, 8)),
			1569 => std_logic_vector(to_unsigned(92, 8)),
			1570 => std_logic_vector(to_unsigned(211, 8)),
			1571 => std_logic_vector(to_unsigned(92, 8)),
			1572 => std_logic_vector(to_unsigned(6, 8)),
			1573 => std_logic_vector(to_unsigned(184, 8)),
			1574 => std_logic_vector(to_unsigned(139, 8)),
			1575 => std_logic_vector(to_unsigned(183, 8)),
			1576 => std_logic_vector(to_unsigned(55, 8)),
			1577 => std_logic_vector(to_unsigned(207, 8)),
			1578 => std_logic_vector(to_unsigned(7, 8)),
			1579 => std_logic_vector(to_unsigned(109, 8)),
			1580 => std_logic_vector(to_unsigned(165, 8)),
			1581 => std_logic_vector(to_unsigned(15, 8)),
			1582 => std_logic_vector(to_unsigned(114, 8)),
			1583 => std_logic_vector(to_unsigned(131, 8)),
			1584 => std_logic_vector(to_unsigned(139, 8)),
			1585 => std_logic_vector(to_unsigned(172, 8)),
			1586 => std_logic_vector(to_unsigned(68, 8)),
			1587 => std_logic_vector(to_unsigned(28, 8)),
			1588 => std_logic_vector(to_unsigned(183, 8)),
			1589 => std_logic_vector(to_unsigned(252, 8)),
			1590 => std_logic_vector(to_unsigned(0, 8)),
			1591 => std_logic_vector(to_unsigned(66, 8)),
			1592 => std_logic_vector(to_unsigned(185, 8)),
			1593 => std_logic_vector(to_unsigned(118, 8)),
			1594 => std_logic_vector(to_unsigned(150, 8)),
			1595 => std_logic_vector(to_unsigned(219, 8)),
			1596 => std_logic_vector(to_unsigned(36, 8)),
			1597 => std_logic_vector(to_unsigned(115, 8)),
			1598 => std_logic_vector(to_unsigned(104, 8)),
			1599 => std_logic_vector(to_unsigned(189, 8)),
			1600 => std_logic_vector(to_unsigned(104, 8)),
			1601 => std_logic_vector(to_unsigned(125, 8)),
			1602 => std_logic_vector(to_unsigned(148, 8)),
			1603 => std_logic_vector(to_unsigned(174, 8)),
			1604 => std_logic_vector(to_unsigned(19, 8)),
			1605 => std_logic_vector(to_unsigned(178, 8)),
			1606 => std_logic_vector(to_unsigned(13, 8)),
			1607 => std_logic_vector(to_unsigned(199, 8)),
			1608 => std_logic_vector(to_unsigned(66, 8)),
			1609 => std_logic_vector(to_unsigned(176, 8)),
			1610 => std_logic_vector(to_unsigned(240, 8)),
			1611 => std_logic_vector(to_unsigned(38, 8)),
			1612 => std_logic_vector(to_unsigned(211, 8)),
			1613 => std_logic_vector(to_unsigned(68, 8)),
			1614 => std_logic_vector(to_unsigned(248, 8)),
			1615 => std_logic_vector(to_unsigned(225, 8)),
			1616 => std_logic_vector(to_unsigned(139, 8)),
			1617 => std_logic_vector(to_unsigned(193, 8)),
			1618 => std_logic_vector(to_unsigned(222, 8)),
			1619 => std_logic_vector(to_unsigned(184, 8)),
			1620 => std_logic_vector(to_unsigned(239, 8)),
			1621 => std_logic_vector(to_unsigned(106, 8)),
			1622 => std_logic_vector(to_unsigned(228, 8)),
			1623 => std_logic_vector(to_unsigned(13, 8)),
			1624 => std_logic_vector(to_unsigned(173, 8)),
			1625 => std_logic_vector(to_unsigned(238, 8)),
			1626 => std_logic_vector(to_unsigned(255, 8)),
			1627 => std_logic_vector(to_unsigned(159, 8)),
			1628 => std_logic_vector(to_unsigned(183, 8)),
			1629 => std_logic_vector(to_unsigned(13, 8)),
			1630 => std_logic_vector(to_unsigned(153, 8)),
			1631 => std_logic_vector(to_unsigned(210, 8)),
			1632 => std_logic_vector(to_unsigned(86, 8)),
			1633 => std_logic_vector(to_unsigned(151, 8)),
			1634 => std_logic_vector(to_unsigned(96, 8)),
			1635 => std_logic_vector(to_unsigned(4, 8)),
			1636 => std_logic_vector(to_unsigned(171, 8)),
			1637 => std_logic_vector(to_unsigned(226, 8)),
			1638 => std_logic_vector(to_unsigned(83, 8)),
			1639 => std_logic_vector(to_unsigned(34, 8)),
			1640 => std_logic_vector(to_unsigned(117, 8)),
			1641 => std_logic_vector(to_unsigned(168, 8)),
			1642 => std_logic_vector(to_unsigned(69, 8)),
			1643 => std_logic_vector(to_unsigned(99, 8)),
			1644 => std_logic_vector(to_unsigned(253, 8)),
			1645 => std_logic_vector(to_unsigned(63, 8)),
			1646 => std_logic_vector(to_unsigned(38, 8)),
			1647 => std_logic_vector(to_unsigned(167, 8)),
			1648 => std_logic_vector(to_unsigned(71, 8)),
			1649 => std_logic_vector(to_unsigned(177, 8)),
			1650 => std_logic_vector(to_unsigned(242, 8)),
			1651 => std_logic_vector(to_unsigned(93, 8)),
			1652 => std_logic_vector(to_unsigned(153, 8)),
			1653 => std_logic_vector(to_unsigned(27, 8)),
			1654 => std_logic_vector(to_unsigned(43, 8)),
			1655 => std_logic_vector(to_unsigned(229, 8)),
			1656 => std_logic_vector(to_unsigned(21, 8)),
			1657 => std_logic_vector(to_unsigned(146, 8)),
			1658 => std_logic_vector(to_unsigned(18, 8)),
			1659 => std_logic_vector(to_unsigned(81, 8)),
			1660 => std_logic_vector(to_unsigned(246, 8)),
			1661 => std_logic_vector(to_unsigned(221, 8)),
			1662 => std_logic_vector(to_unsigned(137, 8)),
			1663 => std_logic_vector(to_unsigned(0, 8)),
			1664 => std_logic_vector(to_unsigned(125, 8)),
			1665 => std_logic_vector(to_unsigned(163, 8)),
			1666 => std_logic_vector(to_unsigned(129, 8)),
			1667 => std_logic_vector(to_unsigned(3, 8)),
			1668 => std_logic_vector(to_unsigned(202, 8)),
			1669 => std_logic_vector(to_unsigned(126, 8)),
			1670 => std_logic_vector(to_unsigned(236, 8)),
			1671 => std_logic_vector(to_unsigned(88, 8)),
			1672 => std_logic_vector(to_unsigned(59, 8)),
			1673 => std_logic_vector(to_unsigned(110, 8)),
			1674 => std_logic_vector(to_unsigned(124, 8)),
			1675 => std_logic_vector(to_unsigned(49, 8)),
			1676 => std_logic_vector(to_unsigned(149, 8)),
			1677 => std_logic_vector(to_unsigned(97, 8)),
			1678 => std_logic_vector(to_unsigned(238, 8)),
			1679 => std_logic_vector(to_unsigned(183, 8)),
			1680 => std_logic_vector(to_unsigned(127, 8)),
			1681 => std_logic_vector(to_unsigned(32, 8)),
			1682 => std_logic_vector(to_unsigned(94, 8)),
			1683 => std_logic_vector(to_unsigned(19, 8)),
			1684 => std_logic_vector(to_unsigned(72, 8)),
			1685 => std_logic_vector(to_unsigned(244, 8)),
			1686 => std_logic_vector(to_unsigned(126, 8)),
			1687 => std_logic_vector(to_unsigned(96, 8)),
			1688 => std_logic_vector(to_unsigned(42, 8)),
			1689 => std_logic_vector(to_unsigned(101, 8)),
			1690 => std_logic_vector(to_unsigned(187, 8)),
			1691 => std_logic_vector(to_unsigned(51, 8)),
			1692 => std_logic_vector(to_unsigned(247, 8)),
			1693 => std_logic_vector(to_unsigned(77, 8)),
			1694 => std_logic_vector(to_unsigned(134, 8)),
			1695 => std_logic_vector(to_unsigned(78, 8)),
			1696 => std_logic_vector(to_unsigned(230, 8)),
			1697 => std_logic_vector(to_unsigned(91, 8)),
			1698 => std_logic_vector(to_unsigned(193, 8)),
			1699 => std_logic_vector(to_unsigned(19, 8)),
			1700 => std_logic_vector(to_unsigned(162, 8)),
			1701 => std_logic_vector(to_unsigned(100, 8)),
			1702 => std_logic_vector(to_unsigned(63, 8)),
			1703 => std_logic_vector(to_unsigned(209, 8)),
			1704 => std_logic_vector(to_unsigned(24, 8)),
			1705 => std_logic_vector(to_unsigned(54, 8)),
			1706 => std_logic_vector(to_unsigned(153, 8)),
			1707 => std_logic_vector(to_unsigned(102, 8)),
			1708 => std_logic_vector(to_unsigned(3, 8)),
			1709 => std_logic_vector(to_unsigned(131, 8)),
			1710 => std_logic_vector(to_unsigned(65, 8)),
			1711 => std_logic_vector(to_unsigned(251, 8)),
			1712 => std_logic_vector(to_unsigned(2, 8)),
			1713 => std_logic_vector(to_unsigned(146, 8)),
			1714 => std_logic_vector(to_unsigned(150, 8)),
			1715 => std_logic_vector(to_unsigned(184, 8)),
			1716 => std_logic_vector(to_unsigned(144, 8)),
			1717 => std_logic_vector(to_unsigned(212, 8)),
			1718 => std_logic_vector(to_unsigned(88, 8)),
			1719 => std_logic_vector(to_unsigned(74, 8)),
			1720 => std_logic_vector(to_unsigned(99, 8)),
			1721 => std_logic_vector(to_unsigned(13, 8)),
			1722 => std_logic_vector(to_unsigned(160, 8)),
			1723 => std_logic_vector(to_unsigned(221, 8)),
			1724 => std_logic_vector(to_unsigned(160, 8)),
			1725 => std_logic_vector(to_unsigned(182, 8)),
			1726 => std_logic_vector(to_unsigned(15, 8)),
			1727 => std_logic_vector(to_unsigned(18, 8)),
			1728 => std_logic_vector(to_unsigned(51, 8)),
			1729 => std_logic_vector(to_unsigned(78, 8)),
			1730 => std_logic_vector(to_unsigned(225, 8)),
			1731 => std_logic_vector(to_unsigned(248, 8)),
			1732 => std_logic_vector(to_unsigned(122, 8)),
			1733 => std_logic_vector(to_unsigned(249, 8)),
			1734 => std_logic_vector(to_unsigned(162, 8)),
			1735 => std_logic_vector(to_unsigned(180, 8)),
			1736 => std_logic_vector(to_unsigned(189, 8)),
			1737 => std_logic_vector(to_unsigned(173, 8)),
			1738 => std_logic_vector(to_unsigned(154, 8)),
			1739 => std_logic_vector(to_unsigned(139, 8)),
			1740 => std_logic_vector(to_unsigned(7, 8)),
			1741 => std_logic_vector(to_unsigned(3, 8)),
			1742 => std_logic_vector(to_unsigned(55, 8)),
			1743 => std_logic_vector(to_unsigned(155, 8)),
			1744 => std_logic_vector(to_unsigned(173, 8)),
			1745 => std_logic_vector(to_unsigned(36, 8)),
			1746 => std_logic_vector(to_unsigned(5, 8)),
			1747 => std_logic_vector(to_unsigned(161, 8)),
			1748 => std_logic_vector(to_unsigned(161, 8)),
			1749 => std_logic_vector(to_unsigned(6, 8)),
			1750 => std_logic_vector(to_unsigned(156, 8)),
			1751 => std_logic_vector(to_unsigned(113, 8)),
			1752 => std_logic_vector(to_unsigned(224, 8)),
			1753 => std_logic_vector(to_unsigned(69, 8)),
			1754 => std_logic_vector(to_unsigned(207, 8)),
			1755 => std_logic_vector(to_unsigned(41, 8)),
			1756 => std_logic_vector(to_unsigned(37, 8)),
			1757 => std_logic_vector(to_unsigned(254, 8)),
			1758 => std_logic_vector(to_unsigned(179, 8)),
			1759 => std_logic_vector(to_unsigned(23, 8)),
			1760 => std_logic_vector(to_unsigned(224, 8)),
			1761 => std_logic_vector(to_unsigned(199, 8)),
			1762 => std_logic_vector(to_unsigned(79, 8)),
			1763 => std_logic_vector(to_unsigned(134, 8)),
			1764 => std_logic_vector(to_unsigned(190, 8)),
			1765 => std_logic_vector(to_unsigned(108, 8)),
			1766 => std_logic_vector(to_unsigned(110, 8)),
			1767 => std_logic_vector(to_unsigned(126, 8)),
			1768 => std_logic_vector(to_unsigned(51, 8)),
			1769 => std_logic_vector(to_unsigned(122, 8)),
			1770 => std_logic_vector(to_unsigned(83, 8)),
			1771 => std_logic_vector(to_unsigned(117, 8)),
			1772 => std_logic_vector(to_unsigned(195, 8)),
			1773 => std_logic_vector(to_unsigned(23, 8)),
			1774 => std_logic_vector(to_unsigned(112, 8)),
			1775 => std_logic_vector(to_unsigned(129, 8)),
			1776 => std_logic_vector(to_unsigned(3, 8)),
			1777 => std_logic_vector(to_unsigned(157, 8)),
			1778 => std_logic_vector(to_unsigned(205, 8)),
			1779 => std_logic_vector(to_unsigned(144, 8)),
			1780 => std_logic_vector(to_unsigned(125, 8)),
			1781 => std_logic_vector(to_unsigned(90, 8)),
			1782 => std_logic_vector(to_unsigned(197, 8)),
			1783 => std_logic_vector(to_unsigned(88, 8)),
			1784 => std_logic_vector(to_unsigned(181, 8)),
			1785 => std_logic_vector(to_unsigned(142, 8)),
			1786 => std_logic_vector(to_unsigned(81, 8)),
			1787 => std_logic_vector(to_unsigned(13, 8)),
			1788 => std_logic_vector(to_unsigned(178, 8)),
			1789 => std_logic_vector(to_unsigned(95, 8)),
			1790 => std_logic_vector(to_unsigned(19, 8)),
			1791 => std_logic_vector(to_unsigned(188, 8)),
			1792 => std_logic_vector(to_unsigned(124, 8)),
			1793 => std_logic_vector(to_unsigned(41, 8)),
			1794 => std_logic_vector(to_unsigned(154, 8)),
			1795 => std_logic_vector(to_unsigned(195, 8)),
			1796 => std_logic_vector(to_unsigned(118, 8)),
			1797 => std_logic_vector(to_unsigned(188, 8)),
			1798 => std_logic_vector(to_unsigned(134, 8)),
			1799 => std_logic_vector(to_unsigned(190, 8)),
			1800 => std_logic_vector(to_unsigned(2, 8)),
			1801 => std_logic_vector(to_unsigned(18, 8)),
			1802 => std_logic_vector(to_unsigned(1, 8)),
			1803 => std_logic_vector(to_unsigned(50, 8)),
			1804 => std_logic_vector(to_unsigned(109, 8)),
			1805 => std_logic_vector(to_unsigned(18, 8)),
			1806 => std_logic_vector(to_unsigned(100, 8)),
			1807 => std_logic_vector(to_unsigned(60, 8)),
			1808 => std_logic_vector(to_unsigned(180, 8)),
			1809 => std_logic_vector(to_unsigned(136, 8)),
			1810 => std_logic_vector(to_unsigned(97, 8)),
			1811 => std_logic_vector(to_unsigned(74, 8)),
			1812 => std_logic_vector(to_unsigned(220, 8)),
			1813 => std_logic_vector(to_unsigned(191, 8)),
			1814 => std_logic_vector(to_unsigned(169, 8)),
			1815 => std_logic_vector(to_unsigned(67, 8)),
			1816 => std_logic_vector(to_unsigned(17, 8)),
			1817 => std_logic_vector(to_unsigned(197, 8)),
			1818 => std_logic_vector(to_unsigned(163, 8)),
			1819 => std_logic_vector(to_unsigned(38, 8)),
			1820 => std_logic_vector(to_unsigned(204, 8)),
			1821 => std_logic_vector(to_unsigned(96, 8)),
			1822 => std_logic_vector(to_unsigned(55, 8)),
			1823 => std_logic_vector(to_unsigned(222, 8)),
			1824 => std_logic_vector(to_unsigned(149, 8)),
			1825 => std_logic_vector(to_unsigned(247, 8)),
			1826 => std_logic_vector(to_unsigned(131, 8)),
			1827 => std_logic_vector(to_unsigned(44, 8)),
			1828 => std_logic_vector(to_unsigned(167, 8)),
			1829 => std_logic_vector(to_unsigned(157, 8)),
			1830 => std_logic_vector(to_unsigned(131, 8)),
			1831 => std_logic_vector(to_unsigned(198, 8)),
			1832 => std_logic_vector(to_unsigned(164, 8)),
			1833 => std_logic_vector(to_unsigned(180, 8)),
			1834 => std_logic_vector(to_unsigned(232, 8)),
			1835 => std_logic_vector(to_unsigned(19, 8)),
			1836 => std_logic_vector(to_unsigned(20, 8)),
			1837 => std_logic_vector(to_unsigned(196, 8)),
			1838 => std_logic_vector(to_unsigned(42, 8)),
			1839 => std_logic_vector(to_unsigned(45, 8)),
			1840 => std_logic_vector(to_unsigned(236, 8)),
			1841 => std_logic_vector(to_unsigned(68, 8)),
			1842 => std_logic_vector(to_unsigned(191, 8)),
			1843 => std_logic_vector(to_unsigned(176, 8)),
			1844 => std_logic_vector(to_unsigned(54, 8)),
			1845 => std_logic_vector(to_unsigned(75, 8)),
			1846 => std_logic_vector(to_unsigned(158, 8)),
			1847 => std_logic_vector(to_unsigned(129, 8)),
			1848 => std_logic_vector(to_unsigned(35, 8)),
			1849 => std_logic_vector(to_unsigned(242, 8)),
			1850 => std_logic_vector(to_unsigned(163, 8)),
			1851 => std_logic_vector(to_unsigned(99, 8)),
			1852 => std_logic_vector(to_unsigned(235, 8)),
			1853 => std_logic_vector(to_unsigned(136, 8)),
			1854 => std_logic_vector(to_unsigned(5, 8)),
			1855 => std_logic_vector(to_unsigned(35, 8)),
			1856 => std_logic_vector(to_unsigned(109, 8)),
			1857 => std_logic_vector(to_unsigned(248, 8)),
			1858 => std_logic_vector(to_unsigned(208, 8)),
			1859 => std_logic_vector(to_unsigned(106, 8)),
			1860 => std_logic_vector(to_unsigned(43, 8)),
			1861 => std_logic_vector(to_unsigned(111, 8)),
			1862 => std_logic_vector(to_unsigned(201, 8)),
			1863 => std_logic_vector(to_unsigned(138, 8)),
			1864 => std_logic_vector(to_unsigned(253, 8)),
			1865 => std_logic_vector(to_unsigned(17, 8)),
			1866 => std_logic_vector(to_unsigned(250, 8)),
			1867 => std_logic_vector(to_unsigned(219, 8)),
			1868 => std_logic_vector(to_unsigned(47, 8)),
			1869 => std_logic_vector(to_unsigned(107, 8)),
			1870 => std_logic_vector(to_unsigned(50, 8)),
			1871 => std_logic_vector(to_unsigned(12, 8)),
			1872 => std_logic_vector(to_unsigned(31, 8)),
			1873 => std_logic_vector(to_unsigned(230, 8)),
			1874 => std_logic_vector(to_unsigned(87, 8)),
			1875 => std_logic_vector(to_unsigned(138, 8)),
			1876 => std_logic_vector(to_unsigned(186, 8)),
			1877 => std_logic_vector(to_unsigned(173, 8)),
			1878 => std_logic_vector(to_unsigned(83, 8)),
			1879 => std_logic_vector(to_unsigned(83, 8)),
			1880 => std_logic_vector(to_unsigned(74, 8)),
			1881 => std_logic_vector(to_unsigned(47, 8)),
			1882 => std_logic_vector(to_unsigned(246, 8)),
			1883 => std_logic_vector(to_unsigned(33, 8)),
			1884 => std_logic_vector(to_unsigned(188, 8)),
			1885 => std_logic_vector(to_unsigned(168, 8)),
			1886 => std_logic_vector(to_unsigned(49, 8)),
			1887 => std_logic_vector(to_unsigned(3, 8)),
			1888 => std_logic_vector(to_unsigned(19, 8)),
			1889 => std_logic_vector(to_unsigned(128, 8)),
			1890 => std_logic_vector(to_unsigned(103, 8)),
			1891 => std_logic_vector(to_unsigned(127, 8)),
			1892 => std_logic_vector(to_unsigned(237, 8)),
			1893 => std_logic_vector(to_unsigned(60, 8)),
			1894 => std_logic_vector(to_unsigned(226, 8)),
			1895 => std_logic_vector(to_unsigned(129, 8)),
			1896 => std_logic_vector(to_unsigned(168, 8)),
			1897 => std_logic_vector(to_unsigned(129, 8)),
			1898 => std_logic_vector(to_unsigned(244, 8)),
			1899 => std_logic_vector(to_unsigned(255, 8)),
			1900 => std_logic_vector(to_unsigned(6, 8)),
			1901 => std_logic_vector(to_unsigned(77, 8)),
			1902 => std_logic_vector(to_unsigned(116, 8)),
			1903 => std_logic_vector(to_unsigned(29, 8)),
			1904 => std_logic_vector(to_unsigned(1, 8)),
			1905 => std_logic_vector(to_unsigned(162, 8)),
			1906 => std_logic_vector(to_unsigned(10, 8)),
			1907 => std_logic_vector(to_unsigned(166, 8)),
			1908 => std_logic_vector(to_unsigned(164, 8)),
			1909 => std_logic_vector(to_unsigned(24, 8)),
			1910 => std_logic_vector(to_unsigned(142, 8)),
			1911 => std_logic_vector(to_unsigned(160, 8)),
			1912 => std_logic_vector(to_unsigned(9, 8)),
			1913 => std_logic_vector(to_unsigned(127, 8)),
			1914 => std_logic_vector(to_unsigned(253, 8)),
			1915 => std_logic_vector(to_unsigned(22, 8)),
			1916 => std_logic_vector(to_unsigned(134, 8)),
			1917 => std_logic_vector(to_unsigned(51, 8)),
			1918 => std_logic_vector(to_unsigned(192, 8)),
			1919 => std_logic_vector(to_unsigned(1, 8)),
			1920 => std_logic_vector(to_unsigned(244, 8)),
			1921 => std_logic_vector(to_unsigned(220, 8)),
			1922 => std_logic_vector(to_unsigned(99, 8)),
			1923 => std_logic_vector(to_unsigned(22, 8)),
			1924 => std_logic_vector(to_unsigned(101, 8)),
			1925 => std_logic_vector(to_unsigned(107, 8)),
			1926 => std_logic_vector(to_unsigned(56, 8)),
			1927 => std_logic_vector(to_unsigned(197, 8)),
			1928 => std_logic_vector(to_unsigned(246, 8)),
			1929 => std_logic_vector(to_unsigned(35, 8)),
			1930 => std_logic_vector(to_unsigned(69, 8)),
			1931 => std_logic_vector(to_unsigned(13, 8)),
			1932 => std_logic_vector(to_unsigned(105, 8)),
			1933 => std_logic_vector(to_unsigned(110, 8)),
			1934 => std_logic_vector(to_unsigned(37, 8)),
			1935 => std_logic_vector(to_unsigned(47, 8)),
			1936 => std_logic_vector(to_unsigned(103, 8)),
			1937 => std_logic_vector(to_unsigned(17, 8)),
			1938 => std_logic_vector(to_unsigned(71, 8)),
			1939 => std_logic_vector(to_unsigned(192, 8)),
			1940 => std_logic_vector(to_unsigned(41, 8)),
			1941 => std_logic_vector(to_unsigned(106, 8)),
			1942 => std_logic_vector(to_unsigned(115, 8)),
			1943 => std_logic_vector(to_unsigned(200, 8)),
			1944 => std_logic_vector(to_unsigned(150, 8)),
			1945 => std_logic_vector(to_unsigned(144, 8)),
			1946 => std_logic_vector(to_unsigned(72, 8)),
			1947 => std_logic_vector(to_unsigned(77, 8)),
			1948 => std_logic_vector(to_unsigned(223, 8)),
			1949 => std_logic_vector(to_unsigned(149, 8)),
			1950 => std_logic_vector(to_unsigned(55, 8)),
			1951 => std_logic_vector(to_unsigned(82, 8)),
			1952 => std_logic_vector(to_unsigned(80, 8)),
			1953 => std_logic_vector(to_unsigned(229, 8)),
			1954 => std_logic_vector(to_unsigned(75, 8)),
			1955 => std_logic_vector(to_unsigned(220, 8)),
			1956 => std_logic_vector(to_unsigned(168, 8)),
			1957 => std_logic_vector(to_unsigned(193, 8)),
			1958 => std_logic_vector(to_unsigned(26, 8)),
			1959 => std_logic_vector(to_unsigned(30, 8)),
			1960 => std_logic_vector(to_unsigned(19, 8)),
			1961 => std_logic_vector(to_unsigned(127, 8)),
			1962 => std_logic_vector(to_unsigned(185, 8)),
			1963 => std_logic_vector(to_unsigned(33, 8)),
			1964 => std_logic_vector(to_unsigned(41, 8)),
			1965 => std_logic_vector(to_unsigned(255, 8)),
			1966 => std_logic_vector(to_unsigned(46, 8)),
			1967 => std_logic_vector(to_unsigned(221, 8)),
			1968 => std_logic_vector(to_unsigned(133, 8)),
			1969 => std_logic_vector(to_unsigned(74, 8)),
			1970 => std_logic_vector(to_unsigned(255, 8)),
			1971 => std_logic_vector(to_unsigned(40, 8)),
			1972 => std_logic_vector(to_unsigned(202, 8)),
			1973 => std_logic_vector(to_unsigned(253, 8)),
			1974 => std_logic_vector(to_unsigned(183, 8)),
			1975 => std_logic_vector(to_unsigned(57, 8)),
			1976 => std_logic_vector(to_unsigned(150, 8)),
			1977 => std_logic_vector(to_unsigned(139, 8)),
			1978 => std_logic_vector(to_unsigned(9, 8)),
			1979 => std_logic_vector(to_unsigned(68, 8)),
			1980 => std_logic_vector(to_unsigned(119, 8)),
			1981 => std_logic_vector(to_unsigned(20, 8)),
			1982 => std_logic_vector(to_unsigned(78, 8)),
			1983 => std_logic_vector(to_unsigned(29, 8)),
			1984 => std_logic_vector(to_unsigned(241, 8)),
			1985 => std_logic_vector(to_unsigned(70, 8)),
			1986 => std_logic_vector(to_unsigned(245, 8)),
			1987 => std_logic_vector(to_unsigned(178, 8)),
			1988 => std_logic_vector(to_unsigned(84, 8)),
			1989 => std_logic_vector(to_unsigned(14, 8)),
			1990 => std_logic_vector(to_unsigned(208, 8)),
			1991 => std_logic_vector(to_unsigned(102, 8)),
			1992 => std_logic_vector(to_unsigned(65, 8)),
			1993 => std_logic_vector(to_unsigned(197, 8)),
			1994 => std_logic_vector(to_unsigned(47, 8)),
			1995 => std_logic_vector(to_unsigned(70, 8)),
			1996 => std_logic_vector(to_unsigned(175, 8)),
			1997 => std_logic_vector(to_unsigned(213, 8)),
			1998 => std_logic_vector(to_unsigned(214, 8)),
			1999 => std_logic_vector(to_unsigned(217, 8)),
			2000 => std_logic_vector(to_unsigned(62, 8)),
			2001 => std_logic_vector(to_unsigned(91, 8)),
			2002 => std_logic_vector(to_unsigned(86, 8)),
			2003 => std_logic_vector(to_unsigned(65, 8)),
			2004 => std_logic_vector(to_unsigned(233, 8)),
			2005 => std_logic_vector(to_unsigned(18, 8)),
			2006 => std_logic_vector(to_unsigned(7, 8)),
			2007 => std_logic_vector(to_unsigned(70, 8)),
			2008 => std_logic_vector(to_unsigned(17, 8)),
			2009 => std_logic_vector(to_unsigned(230, 8)),
			2010 => std_logic_vector(to_unsigned(57, 8)),
			2011 => std_logic_vector(to_unsigned(148, 8)),
			2012 => std_logic_vector(to_unsigned(105, 8)),
			2013 => std_logic_vector(to_unsigned(124, 8)),
			2014 => std_logic_vector(to_unsigned(122, 8)),
			2015 => std_logic_vector(to_unsigned(116, 8)),
			2016 => std_logic_vector(to_unsigned(176, 8)),
			2017 => std_logic_vector(to_unsigned(26, 8)),
			2018 => std_logic_vector(to_unsigned(71, 8)),
			2019 => std_logic_vector(to_unsigned(62, 8)),
			2020 => std_logic_vector(to_unsigned(199, 8)),
			2021 => std_logic_vector(to_unsigned(63, 8)),
			2022 => std_logic_vector(to_unsigned(93, 8)),
			2023 => std_logic_vector(to_unsigned(248, 8)),
			2024 => std_logic_vector(to_unsigned(198, 8)),
			2025 => std_logic_vector(to_unsigned(109, 8)),
			2026 => std_logic_vector(to_unsigned(55, 8)),
			2027 => std_logic_vector(to_unsigned(220, 8)),
			2028 => std_logic_vector(to_unsigned(144, 8)),
			2029 => std_logic_vector(to_unsigned(80, 8)),
			2030 => std_logic_vector(to_unsigned(189, 8)),
			2031 => std_logic_vector(to_unsigned(116, 8)),
			2032 => std_logic_vector(to_unsigned(124, 8)),
			2033 => std_logic_vector(to_unsigned(75, 8)),
			2034 => std_logic_vector(to_unsigned(171, 8)),
			2035 => std_logic_vector(to_unsigned(131, 8)),
			2036 => std_logic_vector(to_unsigned(221, 8)),
			2037 => std_logic_vector(to_unsigned(56, 8)),
			2038 => std_logic_vector(to_unsigned(66, 8)),
			2039 => std_logic_vector(to_unsigned(225, 8)),
			2040 => std_logic_vector(to_unsigned(214, 8)),
			2041 => std_logic_vector(to_unsigned(253, 8)),
			2042 => std_logic_vector(to_unsigned(243, 8)),
			2043 => std_logic_vector(to_unsigned(58, 8)),
			2044 => std_logic_vector(to_unsigned(228, 8)),
			2045 => std_logic_vector(to_unsigned(216, 8)),
			2046 => std_logic_vector(to_unsigned(22, 8)),
			2047 => std_logic_vector(to_unsigned(31, 8)),
			2048 => std_logic_vector(to_unsigned(8, 8)),
			2049 => std_logic_vector(to_unsigned(121, 8)),
			2050 => std_logic_vector(to_unsigned(173, 8)),
			2051 => std_logic_vector(to_unsigned(108, 8)),
			2052 => std_logic_vector(to_unsigned(20, 8)),
			2053 => std_logic_vector(to_unsigned(158, 8)),
			2054 => std_logic_vector(to_unsigned(40, 8)),
			2055 => std_logic_vector(to_unsigned(235, 8)),
			2056 => std_logic_vector(to_unsigned(44, 8)),
			2057 => std_logic_vector(to_unsigned(13, 8)),
			2058 => std_logic_vector(to_unsigned(215, 8)),
			2059 => std_logic_vector(to_unsigned(164, 8)),
			2060 => std_logic_vector(to_unsigned(163, 8)),
			2061 => std_logic_vector(to_unsigned(66, 8)),
			2062 => std_logic_vector(to_unsigned(74, 8)),
			2063 => std_logic_vector(to_unsigned(221, 8)),
			2064 => std_logic_vector(to_unsigned(62, 8)),
			2065 => std_logic_vector(to_unsigned(161, 8)),
			2066 => std_logic_vector(to_unsigned(153, 8)),
			2067 => std_logic_vector(to_unsigned(232, 8)),
			2068 => std_logic_vector(to_unsigned(68, 8)),
			2069 => std_logic_vector(to_unsigned(191, 8)),
			2070 => std_logic_vector(to_unsigned(64, 8)),
			2071 => std_logic_vector(to_unsigned(165, 8)),
			2072 => std_logic_vector(to_unsigned(182, 8)),
			2073 => std_logic_vector(to_unsigned(205, 8)),
			2074 => std_logic_vector(to_unsigned(238, 8)),
			2075 => std_logic_vector(to_unsigned(229, 8)),
			2076 => std_logic_vector(to_unsigned(123, 8)),
			2077 => std_logic_vector(to_unsigned(217, 8)),
			2078 => std_logic_vector(to_unsigned(103, 8)),
			2079 => std_logic_vector(to_unsigned(207, 8)),
			2080 => std_logic_vector(to_unsigned(169, 8)),
			2081 => std_logic_vector(to_unsigned(142, 8)),
			2082 => std_logic_vector(to_unsigned(251, 8)),
			2083 => std_logic_vector(to_unsigned(6, 8)),
			2084 => std_logic_vector(to_unsigned(100, 8)),
			2085 => std_logic_vector(to_unsigned(201, 8)),
			2086 => std_logic_vector(to_unsigned(216, 8)),
			2087 => std_logic_vector(to_unsigned(157, 8)),
			2088 => std_logic_vector(to_unsigned(224, 8)),
			2089 => std_logic_vector(to_unsigned(129, 8)),
			2090 => std_logic_vector(to_unsigned(133, 8)),
			2091 => std_logic_vector(to_unsigned(202, 8)),
			2092 => std_logic_vector(to_unsigned(162, 8)),
			2093 => std_logic_vector(to_unsigned(254, 8)),
			2094 => std_logic_vector(to_unsigned(31, 8)),
			2095 => std_logic_vector(to_unsigned(102, 8)),
			2096 => std_logic_vector(to_unsigned(31, 8)),
			2097 => std_logic_vector(to_unsigned(193, 8)),
			2098 => std_logic_vector(to_unsigned(155, 8)),
			2099 => std_logic_vector(to_unsigned(227, 8)),
			2100 => std_logic_vector(to_unsigned(235, 8)),
			2101 => std_logic_vector(to_unsigned(61, 8)),
			2102 => std_logic_vector(to_unsigned(191, 8)),
			2103 => std_logic_vector(to_unsigned(60, 8)),
			2104 => std_logic_vector(to_unsigned(246, 8)),
			2105 => std_logic_vector(to_unsigned(131, 8)),
			2106 => std_logic_vector(to_unsigned(72, 8)),
			2107 => std_logic_vector(to_unsigned(143, 8)),
			2108 => std_logic_vector(to_unsigned(159, 8)),
			2109 => std_logic_vector(to_unsigned(255, 8)),
			2110 => std_logic_vector(to_unsigned(78, 8)),
			2111 => std_logic_vector(to_unsigned(69, 8)),
			2112 => std_logic_vector(to_unsigned(166, 8)),
			2113 => std_logic_vector(to_unsigned(156, 8)),
			2114 => std_logic_vector(to_unsigned(4, 8)),
			2115 => std_logic_vector(to_unsigned(1, 8)),
			2116 => std_logic_vector(to_unsigned(33, 8)),
			2117 => std_logic_vector(to_unsigned(110, 8)),
			2118 => std_logic_vector(to_unsigned(201, 8)),
			2119 => std_logic_vector(to_unsigned(205, 8)),
			2120 => std_logic_vector(to_unsigned(53, 8)),
			2121 => std_logic_vector(to_unsigned(123, 8)),
			2122 => std_logic_vector(to_unsigned(78, 8)),
			2123 => std_logic_vector(to_unsigned(87, 8)),
			2124 => std_logic_vector(to_unsigned(180, 8)),
			2125 => std_logic_vector(to_unsigned(27, 8)),
			2126 => std_logic_vector(to_unsigned(24, 8)),
			2127 => std_logic_vector(to_unsigned(178, 8)),
			2128 => std_logic_vector(to_unsigned(35, 8)),
			2129 => std_logic_vector(to_unsigned(92, 8)),
			2130 => std_logic_vector(to_unsigned(96, 8)),
			2131 => std_logic_vector(to_unsigned(158, 8)),
			2132 => std_logic_vector(to_unsigned(154, 8)),
			2133 => std_logic_vector(to_unsigned(108, 8)),
			2134 => std_logic_vector(to_unsigned(128, 8)),
			2135 => std_logic_vector(to_unsigned(230, 8)),
			2136 => std_logic_vector(to_unsigned(63, 8)),
			2137 => std_logic_vector(to_unsigned(57, 8)),
			2138 => std_logic_vector(to_unsigned(217, 8)),
			2139 => std_logic_vector(to_unsigned(51, 8)),
			2140 => std_logic_vector(to_unsigned(88, 8)),
			2141 => std_logic_vector(to_unsigned(155, 8)),
			2142 => std_logic_vector(to_unsigned(112, 8)),
			2143 => std_logic_vector(to_unsigned(56, 8)),
			2144 => std_logic_vector(to_unsigned(229, 8)),
			2145 => std_logic_vector(to_unsigned(54, 8)),
			2146 => std_logic_vector(to_unsigned(67, 8)),
			2147 => std_logic_vector(to_unsigned(44, 8)),
			2148 => std_logic_vector(to_unsigned(41, 8)),
			2149 => std_logic_vector(to_unsigned(56, 8)),
			2150 => std_logic_vector(to_unsigned(216, 8)),
			2151 => std_logic_vector(to_unsigned(105, 8)),
			2152 => std_logic_vector(to_unsigned(147, 8)),
			2153 => std_logic_vector(to_unsigned(48, 8)),
			2154 => std_logic_vector(to_unsigned(183, 8)),
			2155 => std_logic_vector(to_unsigned(69, 8)),
			2156 => std_logic_vector(to_unsigned(211, 8)),
			2157 => std_logic_vector(to_unsigned(135, 8)),
			2158 => std_logic_vector(to_unsigned(48, 8)),
			2159 => std_logic_vector(to_unsigned(165, 8)),
			2160 => std_logic_vector(to_unsigned(17, 8)),
			2161 => std_logic_vector(to_unsigned(149, 8)),
			2162 => std_logic_vector(to_unsigned(230, 8)),
			2163 => std_logic_vector(to_unsigned(84, 8)),
			2164 => std_logic_vector(to_unsigned(157, 8)),
			2165 => std_logic_vector(to_unsigned(149, 8)),
			2166 => std_logic_vector(to_unsigned(168, 8)),
			2167 => std_logic_vector(to_unsigned(48, 8)),
			2168 => std_logic_vector(to_unsigned(89, 8)),
			2169 => std_logic_vector(to_unsigned(2, 8)),
			2170 => std_logic_vector(to_unsigned(241, 8)),
			2171 => std_logic_vector(to_unsigned(121, 8)),
			2172 => std_logic_vector(to_unsigned(3, 8)),
			2173 => std_logic_vector(to_unsigned(106, 8)),
			2174 => std_logic_vector(to_unsigned(166, 8)),
			2175 => std_logic_vector(to_unsigned(210, 8)),
			2176 => std_logic_vector(to_unsigned(165, 8)),
			2177 => std_logic_vector(to_unsigned(25, 8)),
			2178 => std_logic_vector(to_unsigned(170, 8)),
			2179 => std_logic_vector(to_unsigned(199, 8)),
			2180 => std_logic_vector(to_unsigned(192, 8)),
			2181 => std_logic_vector(to_unsigned(9, 8)),
			2182 => std_logic_vector(to_unsigned(236, 8)),
			2183 => std_logic_vector(to_unsigned(255, 8)),
			2184 => std_logic_vector(to_unsigned(84, 8)),
			2185 => std_logic_vector(to_unsigned(133, 8)),
			2186 => std_logic_vector(to_unsigned(78, 8)),
			2187 => std_logic_vector(to_unsigned(80, 8)),
			2188 => std_logic_vector(to_unsigned(127, 8)),
			2189 => std_logic_vector(to_unsigned(216, 8)),
			2190 => std_logic_vector(to_unsigned(219, 8)),
			2191 => std_logic_vector(to_unsigned(21, 8)),
			2192 => std_logic_vector(to_unsigned(36, 8)),
			2193 => std_logic_vector(to_unsigned(65, 8)),
			2194 => std_logic_vector(to_unsigned(70, 8)),
			2195 => std_logic_vector(to_unsigned(216, 8)),
			2196 => std_logic_vector(to_unsigned(178, 8)),
			2197 => std_logic_vector(to_unsigned(129, 8)),
			2198 => std_logic_vector(to_unsigned(234, 8)),
			2199 => std_logic_vector(to_unsigned(179, 8)),
			2200 => std_logic_vector(to_unsigned(199, 8)),
			2201 => std_logic_vector(to_unsigned(99, 8)),
			2202 => std_logic_vector(to_unsigned(10, 8)),
			2203 => std_logic_vector(to_unsigned(30, 8)),
			2204 => std_logic_vector(to_unsigned(207, 8)),
			2205 => std_logic_vector(to_unsigned(67, 8)),
			2206 => std_logic_vector(to_unsigned(8, 8)),
			2207 => std_logic_vector(to_unsigned(226, 8)),
			2208 => std_logic_vector(to_unsigned(214, 8)),
			2209 => std_logic_vector(to_unsigned(39, 8)),
			2210 => std_logic_vector(to_unsigned(160, 8)),
			2211 => std_logic_vector(to_unsigned(201, 8)),
			2212 => std_logic_vector(to_unsigned(95, 8)),
			2213 => std_logic_vector(to_unsigned(170, 8)),
			2214 => std_logic_vector(to_unsigned(221, 8)),
			2215 => std_logic_vector(to_unsigned(59, 8)),
			2216 => std_logic_vector(to_unsigned(162, 8)),
			2217 => std_logic_vector(to_unsigned(111, 8)),
			2218 => std_logic_vector(to_unsigned(221, 8)),
			2219 => std_logic_vector(to_unsigned(53, 8)),
			2220 => std_logic_vector(to_unsigned(255, 8)),
			2221 => std_logic_vector(to_unsigned(147, 8)),
			2222 => std_logic_vector(to_unsigned(238, 8)),
			2223 => std_logic_vector(to_unsigned(30, 8)),
			2224 => std_logic_vector(to_unsigned(58, 8)),
			2225 => std_logic_vector(to_unsigned(108, 8)),
			2226 => std_logic_vector(to_unsigned(16, 8)),
			2227 => std_logic_vector(to_unsigned(199, 8)),
			2228 => std_logic_vector(to_unsigned(242, 8)),
			2229 => std_logic_vector(to_unsigned(47, 8)),
			2230 => std_logic_vector(to_unsigned(146, 8)),
			2231 => std_logic_vector(to_unsigned(221, 8)),
			2232 => std_logic_vector(to_unsigned(163, 8)),
			2233 => std_logic_vector(to_unsigned(163, 8)),
			2234 => std_logic_vector(to_unsigned(208, 8)),
			2235 => std_logic_vector(to_unsigned(195, 8)),
			2236 => std_logic_vector(to_unsigned(154, 8)),
			2237 => std_logic_vector(to_unsigned(97, 8)),
			2238 => std_logic_vector(to_unsigned(169, 8)),
			2239 => std_logic_vector(to_unsigned(20, 8)),
			2240 => std_logic_vector(to_unsigned(137, 8)),
			2241 => std_logic_vector(to_unsigned(185, 8)),
			2242 => std_logic_vector(to_unsigned(36, 8)),
			2243 => std_logic_vector(to_unsigned(21, 8)),
			2244 => std_logic_vector(to_unsigned(209, 8)),
			2245 => std_logic_vector(to_unsigned(134, 8)),
			2246 => std_logic_vector(to_unsigned(91, 8)),
			2247 => std_logic_vector(to_unsigned(173, 8)),
			2248 => std_logic_vector(to_unsigned(99, 8)),
			2249 => std_logic_vector(to_unsigned(44, 8)),
			2250 => std_logic_vector(to_unsigned(114, 8)),
			2251 => std_logic_vector(to_unsigned(37, 8)),
			2252 => std_logic_vector(to_unsigned(226, 8)),
			2253 => std_logic_vector(to_unsigned(93, 8)),
			2254 => std_logic_vector(to_unsigned(41, 8)),
			2255 => std_logic_vector(to_unsigned(162, 8)),
			2256 => std_logic_vector(to_unsigned(200, 8)),
			2257 => std_logic_vector(to_unsigned(137, 8)),
			2258 => std_logic_vector(to_unsigned(49, 8)),
			2259 => std_logic_vector(to_unsigned(155, 8)),
			2260 => std_logic_vector(to_unsigned(192, 8)),
			2261 => std_logic_vector(to_unsigned(224, 8)),
			2262 => std_logic_vector(to_unsigned(244, 8)),
			2263 => std_logic_vector(to_unsigned(255, 8)),
			2264 => std_logic_vector(to_unsigned(47, 8)),
			2265 => std_logic_vector(to_unsigned(54, 8)),
			2266 => std_logic_vector(to_unsigned(112, 8)),
			2267 => std_logic_vector(to_unsigned(118, 8)),
			2268 => std_logic_vector(to_unsigned(42, 8)),
			2269 => std_logic_vector(to_unsigned(40, 8)),
			2270 => std_logic_vector(to_unsigned(154, 8)),
			2271 => std_logic_vector(to_unsigned(174, 8)),
			2272 => std_logic_vector(to_unsigned(240, 8)),
			2273 => std_logic_vector(to_unsigned(199, 8)),
			2274 => std_logic_vector(to_unsigned(246, 8)),
			2275 => std_logic_vector(to_unsigned(109, 8)),
			2276 => std_logic_vector(to_unsigned(84, 8)),
			2277 => std_logic_vector(to_unsigned(196, 8)),
			2278 => std_logic_vector(to_unsigned(41, 8)),
			2279 => std_logic_vector(to_unsigned(68, 8)),
			2280 => std_logic_vector(to_unsigned(82, 8)),
			2281 => std_logic_vector(to_unsigned(40, 8)),
			2282 => std_logic_vector(to_unsigned(154, 8)),
			2283 => std_logic_vector(to_unsigned(13, 8)),
			2284 => std_logic_vector(to_unsigned(57, 8)),
			2285 => std_logic_vector(to_unsigned(129, 8)),
			2286 => std_logic_vector(to_unsigned(9, 8)),
			2287 => std_logic_vector(to_unsigned(160, 8)),
			2288 => std_logic_vector(to_unsigned(230, 8)),
			2289 => std_logic_vector(to_unsigned(190, 8)),
			2290 => std_logic_vector(to_unsigned(136, 8)),
			2291 => std_logic_vector(to_unsigned(115, 8)),
			2292 => std_logic_vector(to_unsigned(233, 8)),
			2293 => std_logic_vector(to_unsigned(203, 8)),
			2294 => std_logic_vector(to_unsigned(213, 8)),
			2295 => std_logic_vector(to_unsigned(244, 8)),
			2296 => std_logic_vector(to_unsigned(22, 8)),
			2297 => std_logic_vector(to_unsigned(156, 8)),
			2298 => std_logic_vector(to_unsigned(59, 8)),
			2299 => std_logic_vector(to_unsigned(178, 8)),
			2300 => std_logic_vector(to_unsigned(135, 8)),
			2301 => std_logic_vector(to_unsigned(242, 8)),
			2302 => std_logic_vector(to_unsigned(5, 8)),
			2303 => std_logic_vector(to_unsigned(195, 8)),
			2304 => std_logic_vector(to_unsigned(237, 8)),
			2305 => std_logic_vector(to_unsigned(110, 8)),
			2306 => std_logic_vector(to_unsigned(38, 8)),
			2307 => std_logic_vector(to_unsigned(44, 8)),
			2308 => std_logic_vector(to_unsigned(123, 8)),
			2309 => std_logic_vector(to_unsigned(58, 8)),
			2310 => std_logic_vector(to_unsigned(34, 8)),
			2311 => std_logic_vector(to_unsigned(73, 8)),
			2312 => std_logic_vector(to_unsigned(47, 8)),
			2313 => std_logic_vector(to_unsigned(20, 8)),
			2314 => std_logic_vector(to_unsigned(162, 8)),
			2315 => std_logic_vector(to_unsigned(94, 8)),
			2316 => std_logic_vector(to_unsigned(81, 8)),
			2317 => std_logic_vector(to_unsigned(7, 8)),
			2318 => std_logic_vector(to_unsigned(60, 8)),
			2319 => std_logic_vector(to_unsigned(198, 8)),
			2320 => std_logic_vector(to_unsigned(161, 8)),
			2321 => std_logic_vector(to_unsigned(208, 8)),
			2322 => std_logic_vector(to_unsigned(121, 8)),
			2323 => std_logic_vector(to_unsigned(103, 8)),
			2324 => std_logic_vector(to_unsigned(178, 8)),
			2325 => std_logic_vector(to_unsigned(20, 8)),
			2326 => std_logic_vector(to_unsigned(37, 8)),
			2327 => std_logic_vector(to_unsigned(49, 8)),
			2328 => std_logic_vector(to_unsigned(178, 8)),
			2329 => std_logic_vector(to_unsigned(91, 8)),
			2330 => std_logic_vector(to_unsigned(167, 8)),
			2331 => std_logic_vector(to_unsigned(32, 8)),
			2332 => std_logic_vector(to_unsigned(182, 8)),
			2333 => std_logic_vector(to_unsigned(28, 8)),
			2334 => std_logic_vector(to_unsigned(149, 8)),
			2335 => std_logic_vector(to_unsigned(167, 8)),
			2336 => std_logic_vector(to_unsigned(98, 8)),
			2337 => std_logic_vector(to_unsigned(83, 8)),
			2338 => std_logic_vector(to_unsigned(43, 8)),
			2339 => std_logic_vector(to_unsigned(5, 8)),
			2340 => std_logic_vector(to_unsigned(180, 8)),
			2341 => std_logic_vector(to_unsigned(94, 8)),
			2342 => std_logic_vector(to_unsigned(69, 8)),
			2343 => std_logic_vector(to_unsigned(177, 8)),
			2344 => std_logic_vector(to_unsigned(99, 8)),
			2345 => std_logic_vector(to_unsigned(83, 8)),
			2346 => std_logic_vector(to_unsigned(26, 8)),
			2347 => std_logic_vector(to_unsigned(3, 8)),
			2348 => std_logic_vector(to_unsigned(234, 8)),
			2349 => std_logic_vector(to_unsigned(231, 8)),
			2350 => std_logic_vector(to_unsigned(45, 8)),
			2351 => std_logic_vector(to_unsigned(144, 8)),
			2352 => std_logic_vector(to_unsigned(112, 8)),
			2353 => std_logic_vector(to_unsigned(214, 8)),
			2354 => std_logic_vector(to_unsigned(208, 8)),
			2355 => std_logic_vector(to_unsigned(179, 8)),
			2356 => std_logic_vector(to_unsigned(36, 8)),
			2357 => std_logic_vector(to_unsigned(72, 8)),
			2358 => std_logic_vector(to_unsigned(186, 8)),
			2359 => std_logic_vector(to_unsigned(62, 8)),
			2360 => std_logic_vector(to_unsigned(7, 8)),
			2361 => std_logic_vector(to_unsigned(61, 8)),
			2362 => std_logic_vector(to_unsigned(39, 8)),
			2363 => std_logic_vector(to_unsigned(117, 8)),
			2364 => std_logic_vector(to_unsigned(107, 8)),
			2365 => std_logic_vector(to_unsigned(252, 8)),
			2366 => std_logic_vector(to_unsigned(138, 8)),
			2367 => std_logic_vector(to_unsigned(149, 8)),
			2368 => std_logic_vector(to_unsigned(57, 8)),
			2369 => std_logic_vector(to_unsigned(76, 8)),
			2370 => std_logic_vector(to_unsigned(135, 8)),
			2371 => std_logic_vector(to_unsigned(201, 8)),
			2372 => std_logic_vector(to_unsigned(46, 8)),
			2373 => std_logic_vector(to_unsigned(58, 8)),
			2374 => std_logic_vector(to_unsigned(104, 8)),
			2375 => std_logic_vector(to_unsigned(12, 8)),
			2376 => std_logic_vector(to_unsigned(84, 8)),
			2377 => std_logic_vector(to_unsigned(103, 8)),
			2378 => std_logic_vector(to_unsigned(83, 8)),
			2379 => std_logic_vector(to_unsigned(121, 8)),
			2380 => std_logic_vector(to_unsigned(229, 8)),
			2381 => std_logic_vector(to_unsigned(235, 8)),
			2382 => std_logic_vector(to_unsigned(208, 8)),
			2383 => std_logic_vector(to_unsigned(219, 8)),
			2384 => std_logic_vector(to_unsigned(171, 8)),
			2385 => std_logic_vector(to_unsigned(181, 8)),
			2386 => std_logic_vector(to_unsigned(171, 8)),
			2387 => std_logic_vector(to_unsigned(187, 8)),
			2388 => std_logic_vector(to_unsigned(184, 8)),
			2389 => std_logic_vector(to_unsigned(22, 8)),
			2390 => std_logic_vector(to_unsigned(215, 8)),
			2391 => std_logic_vector(to_unsigned(64, 8)),
			2392 => std_logic_vector(to_unsigned(55, 8)),
			2393 => std_logic_vector(to_unsigned(111, 8)),
			2394 => std_logic_vector(to_unsigned(122, 8)),
			2395 => std_logic_vector(to_unsigned(19, 8)),
			2396 => std_logic_vector(to_unsigned(141, 8)),
			2397 => std_logic_vector(to_unsigned(135, 8)),
			2398 => std_logic_vector(to_unsigned(178, 8)),
			2399 => std_logic_vector(to_unsigned(150, 8)),
			2400 => std_logic_vector(to_unsigned(244, 8)),
			2401 => std_logic_vector(to_unsigned(135, 8)),
			2402 => std_logic_vector(to_unsigned(70, 8)),
			2403 => std_logic_vector(to_unsigned(43, 8)),
			2404 => std_logic_vector(to_unsigned(51, 8)),
			2405 => std_logic_vector(to_unsigned(57, 8)),
			2406 => std_logic_vector(to_unsigned(31, 8)),
			2407 => std_logic_vector(to_unsigned(99, 8)),
			2408 => std_logic_vector(to_unsigned(63, 8)),
			2409 => std_logic_vector(to_unsigned(237, 8)),
			2410 => std_logic_vector(to_unsigned(167, 8)),
			2411 => std_logic_vector(to_unsigned(155, 8)),
			2412 => std_logic_vector(to_unsigned(229, 8)),
			2413 => std_logic_vector(to_unsigned(51, 8)),
			2414 => std_logic_vector(to_unsigned(245, 8)),
			2415 => std_logic_vector(to_unsigned(163, 8)),
			2416 => std_logic_vector(to_unsigned(109, 8)),
			2417 => std_logic_vector(to_unsigned(239, 8)),
			2418 => std_logic_vector(to_unsigned(172, 8)),
			2419 => std_logic_vector(to_unsigned(52, 8)),
			2420 => std_logic_vector(to_unsigned(91, 8)),
			2421 => std_logic_vector(to_unsigned(200, 8)),
			2422 => std_logic_vector(to_unsigned(118, 8)),
			2423 => std_logic_vector(to_unsigned(66, 8)),
			2424 => std_logic_vector(to_unsigned(4, 8)),
			2425 => std_logic_vector(to_unsigned(182, 8)),
			2426 => std_logic_vector(to_unsigned(52, 8)),
			2427 => std_logic_vector(to_unsigned(74, 8)),
			2428 => std_logic_vector(to_unsigned(140, 8)),
			2429 => std_logic_vector(to_unsigned(33, 8)),
			2430 => std_logic_vector(to_unsigned(207, 8)),
			2431 => std_logic_vector(to_unsigned(74, 8)),
			2432 => std_logic_vector(to_unsigned(105, 8)),
			2433 => std_logic_vector(to_unsigned(66, 8)),
			2434 => std_logic_vector(to_unsigned(82, 8)),
			2435 => std_logic_vector(to_unsigned(151, 8)),
			2436 => std_logic_vector(to_unsigned(197, 8)),
			2437 => std_logic_vector(to_unsigned(4, 8)),
			2438 => std_logic_vector(to_unsigned(215, 8)),
			2439 => std_logic_vector(to_unsigned(218, 8)),
			2440 => std_logic_vector(to_unsigned(150, 8)),
			2441 => std_logic_vector(to_unsigned(22, 8)),
			2442 => std_logic_vector(to_unsigned(28, 8)),
			2443 => std_logic_vector(to_unsigned(145, 8)),
			2444 => std_logic_vector(to_unsigned(27, 8)),
			2445 => std_logic_vector(to_unsigned(44, 8)),
			2446 => std_logic_vector(to_unsigned(216, 8)),
			2447 => std_logic_vector(to_unsigned(112, 8)),
			2448 => std_logic_vector(to_unsigned(218, 8)),
			2449 => std_logic_vector(to_unsigned(220, 8)),
			2450 => std_logic_vector(to_unsigned(182, 8)),
			2451 => std_logic_vector(to_unsigned(191, 8)),
			2452 => std_logic_vector(to_unsigned(10, 8)),
			2453 => std_logic_vector(to_unsigned(2, 8)),
			2454 => std_logic_vector(to_unsigned(158, 8)),
			2455 => std_logic_vector(to_unsigned(82, 8)),
			2456 => std_logic_vector(to_unsigned(199, 8)),
			2457 => std_logic_vector(to_unsigned(97, 8)),
			2458 => std_logic_vector(to_unsigned(150, 8)),
			2459 => std_logic_vector(to_unsigned(168, 8)),
			2460 => std_logic_vector(to_unsigned(231, 8)),
			2461 => std_logic_vector(to_unsigned(244, 8)),
			2462 => std_logic_vector(to_unsigned(216, 8)),
			2463 => std_logic_vector(to_unsigned(4, 8)),
			2464 => std_logic_vector(to_unsigned(171, 8)),
			2465 => std_logic_vector(to_unsigned(108, 8)),
			2466 => std_logic_vector(to_unsigned(224, 8)),
			2467 => std_logic_vector(to_unsigned(92, 8)),
			2468 => std_logic_vector(to_unsigned(190, 8)),
			2469 => std_logic_vector(to_unsigned(252, 8)),
			2470 => std_logic_vector(to_unsigned(197, 8)),
			2471 => std_logic_vector(to_unsigned(202, 8)),
			2472 => std_logic_vector(to_unsigned(244, 8)),
			2473 => std_logic_vector(to_unsigned(7, 8)),
			2474 => std_logic_vector(to_unsigned(187, 8)),
			2475 => std_logic_vector(to_unsigned(28, 8)),
			2476 => std_logic_vector(to_unsigned(102, 8)),
			2477 => std_logic_vector(to_unsigned(43, 8)),
			2478 => std_logic_vector(to_unsigned(33, 8)),
			2479 => std_logic_vector(to_unsigned(191, 8)),
			2480 => std_logic_vector(to_unsigned(21, 8)),
			2481 => std_logic_vector(to_unsigned(15, 8)),
			2482 => std_logic_vector(to_unsigned(226, 8)),
			2483 => std_logic_vector(to_unsigned(204, 8)),
			2484 => std_logic_vector(to_unsigned(252, 8)),
			2485 => std_logic_vector(to_unsigned(224, 8)),
			2486 => std_logic_vector(to_unsigned(217, 8)),
			2487 => std_logic_vector(to_unsigned(110, 8)),
			2488 => std_logic_vector(to_unsigned(75, 8)),
			2489 => std_logic_vector(to_unsigned(146, 8)),
			2490 => std_logic_vector(to_unsigned(51, 8)),
			2491 => std_logic_vector(to_unsigned(50, 8)),
			2492 => std_logic_vector(to_unsigned(130, 8)),
			2493 => std_logic_vector(to_unsigned(210, 8)),
			2494 => std_logic_vector(to_unsigned(48, 8)),
			2495 => std_logic_vector(to_unsigned(41, 8)),
			2496 => std_logic_vector(to_unsigned(78, 8)),
			2497 => std_logic_vector(to_unsigned(253, 8)),
			2498 => std_logic_vector(to_unsigned(133, 8)),
			2499 => std_logic_vector(to_unsigned(239, 8)),
			2500 => std_logic_vector(to_unsigned(67, 8)),
			2501 => std_logic_vector(to_unsigned(72, 8)),
			2502 => std_logic_vector(to_unsigned(93, 8)),
			2503 => std_logic_vector(to_unsigned(96, 8)),
			2504 => std_logic_vector(to_unsigned(94, 8)),
			2505 => std_logic_vector(to_unsigned(147, 8)),
			2506 => std_logic_vector(to_unsigned(112, 8)),
			2507 => std_logic_vector(to_unsigned(33, 8)),
			2508 => std_logic_vector(to_unsigned(195, 8)),
			2509 => std_logic_vector(to_unsigned(186, 8)),
			2510 => std_logic_vector(to_unsigned(204, 8)),
			2511 => std_logic_vector(to_unsigned(106, 8)),
			2512 => std_logic_vector(to_unsigned(90, 8)),
			2513 => std_logic_vector(to_unsigned(230, 8)),
			2514 => std_logic_vector(to_unsigned(47, 8)),
			2515 => std_logic_vector(to_unsigned(52, 8)),
			2516 => std_logic_vector(to_unsigned(67, 8)),
			2517 => std_logic_vector(to_unsigned(133, 8)),
			2518 => std_logic_vector(to_unsigned(149, 8)),
			2519 => std_logic_vector(to_unsigned(50, 8)),
			2520 => std_logic_vector(to_unsigned(53, 8)),
			2521 => std_logic_vector(to_unsigned(23, 8)),
			2522 => std_logic_vector(to_unsigned(52, 8)),
			2523 => std_logic_vector(to_unsigned(22, 8)),
			2524 => std_logic_vector(to_unsigned(220, 8)),
			2525 => std_logic_vector(to_unsigned(93, 8)),
			2526 => std_logic_vector(to_unsigned(41, 8)),
			2527 => std_logic_vector(to_unsigned(90, 8)),
			2528 => std_logic_vector(to_unsigned(30, 8)),
			2529 => std_logic_vector(to_unsigned(23, 8)),
			2530 => std_logic_vector(to_unsigned(217, 8)),
			2531 => std_logic_vector(to_unsigned(47, 8)),
			2532 => std_logic_vector(to_unsigned(225, 8)),
			2533 => std_logic_vector(to_unsigned(1, 8)),
			2534 => std_logic_vector(to_unsigned(220, 8)),
			2535 => std_logic_vector(to_unsigned(49, 8)),
			2536 => std_logic_vector(to_unsigned(118, 8)),
			2537 => std_logic_vector(to_unsigned(53, 8)),
			2538 => std_logic_vector(to_unsigned(144, 8)),
			2539 => std_logic_vector(to_unsigned(160, 8)),
			2540 => std_logic_vector(to_unsigned(211, 8)),
			2541 => std_logic_vector(to_unsigned(36, 8)),
			2542 => std_logic_vector(to_unsigned(47, 8)),
			2543 => std_logic_vector(to_unsigned(113, 8)),
			2544 => std_logic_vector(to_unsigned(111, 8)),
			2545 => std_logic_vector(to_unsigned(76, 8)),
			2546 => std_logic_vector(to_unsigned(144, 8)),
			2547 => std_logic_vector(to_unsigned(12, 8)),
			2548 => std_logic_vector(to_unsigned(195, 8)),
			2549 => std_logic_vector(to_unsigned(144, 8)),
			2550 => std_logic_vector(to_unsigned(58, 8)),
			2551 => std_logic_vector(to_unsigned(212, 8)),
			2552 => std_logic_vector(to_unsigned(195, 8)),
			2553 => std_logic_vector(to_unsigned(30, 8)),
			2554 => std_logic_vector(to_unsigned(114, 8)),
			2555 => std_logic_vector(to_unsigned(128, 8)),
			2556 => std_logic_vector(to_unsigned(49, 8)),
			2557 => std_logic_vector(to_unsigned(40, 8)),
			2558 => std_logic_vector(to_unsigned(51, 8)),
			2559 => std_logic_vector(to_unsigned(224, 8)),
			2560 => std_logic_vector(to_unsigned(233, 8)),
			2561 => std_logic_vector(to_unsigned(33, 8)),
			2562 => std_logic_vector(to_unsigned(56, 8)),
			2563 => std_logic_vector(to_unsigned(79, 8)),
			2564 => std_logic_vector(to_unsigned(126, 8)),
			2565 => std_logic_vector(to_unsigned(46, 8)),
			2566 => std_logic_vector(to_unsigned(80, 8)),
			2567 => std_logic_vector(to_unsigned(99, 8)),
			2568 => std_logic_vector(to_unsigned(72, 8)),
			2569 => std_logic_vector(to_unsigned(255, 8)),
			2570 => std_logic_vector(to_unsigned(222, 8)),
			2571 => std_logic_vector(to_unsigned(244, 8)),
			2572 => std_logic_vector(to_unsigned(243, 8)),
			2573 => std_logic_vector(to_unsigned(0, 8)),
			2574 => std_logic_vector(to_unsigned(224, 8)),
			2575 => std_logic_vector(to_unsigned(149, 8)),
			2576 => std_logic_vector(to_unsigned(234, 8)),
			2577 => std_logic_vector(to_unsigned(42, 8)),
			2578 => std_logic_vector(to_unsigned(188, 8)),
			2579 => std_logic_vector(to_unsigned(31, 8)),
			2580 => std_logic_vector(to_unsigned(107, 8)),
			2581 => std_logic_vector(to_unsigned(27, 8)),
			2582 => std_logic_vector(to_unsigned(199, 8)),
			2583 => std_logic_vector(to_unsigned(50, 8)),
			2584 => std_logic_vector(to_unsigned(195, 8)),
			2585 => std_logic_vector(to_unsigned(169, 8)),
			2586 => std_logic_vector(to_unsigned(193, 8)),
			2587 => std_logic_vector(to_unsigned(26, 8)),
			2588 => std_logic_vector(to_unsigned(153, 8)),
			2589 => std_logic_vector(to_unsigned(18, 8)),
			2590 => std_logic_vector(to_unsigned(10, 8)),
			2591 => std_logic_vector(to_unsigned(162, 8)),
			2592 => std_logic_vector(to_unsigned(123, 8)),
			2593 => std_logic_vector(to_unsigned(34, 8)),
			2594 => std_logic_vector(to_unsigned(251, 8)),
			2595 => std_logic_vector(to_unsigned(134, 8)),
			2596 => std_logic_vector(to_unsigned(99, 8)),
			2597 => std_logic_vector(to_unsigned(232, 8)),
			2598 => std_logic_vector(to_unsigned(6, 8)),
			2599 => std_logic_vector(to_unsigned(225, 8)),
			2600 => std_logic_vector(to_unsigned(180, 8)),
			2601 => std_logic_vector(to_unsigned(56, 8)),
			2602 => std_logic_vector(to_unsigned(205, 8)),
			2603 => std_logic_vector(to_unsigned(127, 8)),
			2604 => std_logic_vector(to_unsigned(33, 8)),
			2605 => std_logic_vector(to_unsigned(41, 8)),
			2606 => std_logic_vector(to_unsigned(83, 8)),
			2607 => std_logic_vector(to_unsigned(245, 8)),
			2608 => std_logic_vector(to_unsigned(144, 8)),
			2609 => std_logic_vector(to_unsigned(190, 8)),
			2610 => std_logic_vector(to_unsigned(193, 8)),
			2611 => std_logic_vector(to_unsigned(37, 8)),
			2612 => std_logic_vector(to_unsigned(149, 8)),
			2613 => std_logic_vector(to_unsigned(217, 8)),
			2614 => std_logic_vector(to_unsigned(42, 8)),
			2615 => std_logic_vector(to_unsigned(192, 8)),
			2616 => std_logic_vector(to_unsigned(183, 8)),
			2617 => std_logic_vector(to_unsigned(250, 8)),
			2618 => std_logic_vector(to_unsigned(109, 8)),
			2619 => std_logic_vector(to_unsigned(221, 8)),
			2620 => std_logic_vector(to_unsigned(112, 8)),
			2621 => std_logic_vector(to_unsigned(215, 8)),
			2622 => std_logic_vector(to_unsigned(183, 8)),
			2623 => std_logic_vector(to_unsigned(122, 8)),
			2624 => std_logic_vector(to_unsigned(114, 8)),
			2625 => std_logic_vector(to_unsigned(213, 8)),
			2626 => std_logic_vector(to_unsigned(26, 8)),
			2627 => std_logic_vector(to_unsigned(40, 8)),
			2628 => std_logic_vector(to_unsigned(216, 8)),
			2629 => std_logic_vector(to_unsigned(222, 8)),
			2630 => std_logic_vector(to_unsigned(248, 8)),
			2631 => std_logic_vector(to_unsigned(142, 8)),
			2632 => std_logic_vector(to_unsigned(25, 8)),
			2633 => std_logic_vector(to_unsigned(175, 8)),
			2634 => std_logic_vector(to_unsigned(247, 8)),
			2635 => std_logic_vector(to_unsigned(32, 8)),
			2636 => std_logic_vector(to_unsigned(185, 8)),
			2637 => std_logic_vector(to_unsigned(56, 8)),
			2638 => std_logic_vector(to_unsigned(50, 8)),
			2639 => std_logic_vector(to_unsigned(118, 8)),
			2640 => std_logic_vector(to_unsigned(254, 8)),
			2641 => std_logic_vector(to_unsigned(58, 8)),
			2642 => std_logic_vector(to_unsigned(215, 8)),
			2643 => std_logic_vector(to_unsigned(235, 8)),
			2644 => std_logic_vector(to_unsigned(51, 8)),
			2645 => std_logic_vector(to_unsigned(9, 8)),
			2646 => std_logic_vector(to_unsigned(90, 8)),
			2647 => std_logic_vector(to_unsigned(21, 8)),
			2648 => std_logic_vector(to_unsigned(68, 8)),
			2649 => std_logic_vector(to_unsigned(231, 8)),
			2650 => std_logic_vector(to_unsigned(206, 8)),
			2651 => std_logic_vector(to_unsigned(88, 8)),
			2652 => std_logic_vector(to_unsigned(63, 8)),
			2653 => std_logic_vector(to_unsigned(38, 8)),
			2654 => std_logic_vector(to_unsigned(132, 8)),
			2655 => std_logic_vector(to_unsigned(220, 8)),
			2656 => std_logic_vector(to_unsigned(34, 8)),
			2657 => std_logic_vector(to_unsigned(75, 8)),
			2658 => std_logic_vector(to_unsigned(200, 8)),
			2659 => std_logic_vector(to_unsigned(248, 8)),
			2660 => std_logic_vector(to_unsigned(188, 8)),
			2661 => std_logic_vector(to_unsigned(169, 8)),
			2662 => std_logic_vector(to_unsigned(100, 8)),
			2663 => std_logic_vector(to_unsigned(235, 8)),
			2664 => std_logic_vector(to_unsigned(112, 8)),
			2665 => std_logic_vector(to_unsigned(70, 8)),
			2666 => std_logic_vector(to_unsigned(122, 8)),
			2667 => std_logic_vector(to_unsigned(11, 8)),
			2668 => std_logic_vector(to_unsigned(137, 8)),
			2669 => std_logic_vector(to_unsigned(151, 8)),
			2670 => std_logic_vector(to_unsigned(211, 8)),
			2671 => std_logic_vector(to_unsigned(5, 8)),
			2672 => std_logic_vector(to_unsigned(200, 8)),
			2673 => std_logic_vector(to_unsigned(151, 8)),
			2674 => std_logic_vector(to_unsigned(192, 8)),
			2675 => std_logic_vector(to_unsigned(124, 8)),
			2676 => std_logic_vector(to_unsigned(26, 8)),
			2677 => std_logic_vector(to_unsigned(182, 8)),
			2678 => std_logic_vector(to_unsigned(48, 8)),
			2679 => std_logic_vector(to_unsigned(183, 8)),
			2680 => std_logic_vector(to_unsigned(240, 8)),
			2681 => std_logic_vector(to_unsigned(111, 8)),
			2682 => std_logic_vector(to_unsigned(22, 8)),
			2683 => std_logic_vector(to_unsigned(236, 8)),
			2684 => std_logic_vector(to_unsigned(214, 8)),
			2685 => std_logic_vector(to_unsigned(119, 8)),
			2686 => std_logic_vector(to_unsigned(197, 8)),
			2687 => std_logic_vector(to_unsigned(73, 8)),
			2688 => std_logic_vector(to_unsigned(57, 8)),
			2689 => std_logic_vector(to_unsigned(224, 8)),
			2690 => std_logic_vector(to_unsigned(213, 8)),
			2691 => std_logic_vector(to_unsigned(190, 8)),
			2692 => std_logic_vector(to_unsigned(67, 8)),
			2693 => std_logic_vector(to_unsigned(193, 8)),
			2694 => std_logic_vector(to_unsigned(18, 8)),
			2695 => std_logic_vector(to_unsigned(195, 8)),
			2696 => std_logic_vector(to_unsigned(75, 8)),
			2697 => std_logic_vector(to_unsigned(44, 8)),
			2698 => std_logic_vector(to_unsigned(234, 8)),
			2699 => std_logic_vector(to_unsigned(146, 8)),
			2700 => std_logic_vector(to_unsigned(74, 8)),
			2701 => std_logic_vector(to_unsigned(83, 8)),
			2702 => std_logic_vector(to_unsigned(178, 8)),
			2703 => std_logic_vector(to_unsigned(215, 8)),
			2704 => std_logic_vector(to_unsigned(82, 8)),
			2705 => std_logic_vector(to_unsigned(114, 8)),
			2706 => std_logic_vector(to_unsigned(98, 8)),
			2707 => std_logic_vector(to_unsigned(25, 8)),
			2708 => std_logic_vector(to_unsigned(15, 8)),
			2709 => std_logic_vector(to_unsigned(243, 8)),
			2710 => std_logic_vector(to_unsigned(114, 8)),
			2711 => std_logic_vector(to_unsigned(153, 8)),
			2712 => std_logic_vector(to_unsigned(186, 8)),
			2713 => std_logic_vector(to_unsigned(217, 8)),
			2714 => std_logic_vector(to_unsigned(251, 8)),
			2715 => std_logic_vector(to_unsigned(121, 8)),
			2716 => std_logic_vector(to_unsigned(135, 8)),
			2717 => std_logic_vector(to_unsigned(52, 8)),
			2718 => std_logic_vector(to_unsigned(236, 8)),
			2719 => std_logic_vector(to_unsigned(43, 8)),
			2720 => std_logic_vector(to_unsigned(24, 8)),
			2721 => std_logic_vector(to_unsigned(67, 8)),
			2722 => std_logic_vector(to_unsigned(91, 8)),
			2723 => std_logic_vector(to_unsigned(153, 8)),
			2724 => std_logic_vector(to_unsigned(22, 8)),
			2725 => std_logic_vector(to_unsigned(83, 8)),
			2726 => std_logic_vector(to_unsigned(172, 8)),
			2727 => std_logic_vector(to_unsigned(251, 8)),
			2728 => std_logic_vector(to_unsigned(180, 8)),
			2729 => std_logic_vector(to_unsigned(229, 8)),
			2730 => std_logic_vector(to_unsigned(81, 8)),
			2731 => std_logic_vector(to_unsigned(196, 8)),
			2732 => std_logic_vector(to_unsigned(202, 8)),
			2733 => std_logic_vector(to_unsigned(125, 8)),
			2734 => std_logic_vector(to_unsigned(193, 8)),
			2735 => std_logic_vector(to_unsigned(111, 8)),
			2736 => std_logic_vector(to_unsigned(59, 8)),
			2737 => std_logic_vector(to_unsigned(48, 8)),
			2738 => std_logic_vector(to_unsigned(30, 8)),
			2739 => std_logic_vector(to_unsigned(213, 8)),
			2740 => std_logic_vector(to_unsigned(15, 8)),
			2741 => std_logic_vector(to_unsigned(216, 8)),
			2742 => std_logic_vector(to_unsigned(199, 8)),
			2743 => std_logic_vector(to_unsigned(53, 8)),
			2744 => std_logic_vector(to_unsigned(114, 8)),
			2745 => std_logic_vector(to_unsigned(133, 8)),
			2746 => std_logic_vector(to_unsigned(200, 8)),
			2747 => std_logic_vector(to_unsigned(129, 8)),
			2748 => std_logic_vector(to_unsigned(85, 8)),
			2749 => std_logic_vector(to_unsigned(102, 8)),
			2750 => std_logic_vector(to_unsigned(221, 8)),
			2751 => std_logic_vector(to_unsigned(62, 8)),
			2752 => std_logic_vector(to_unsigned(63, 8)),
			2753 => std_logic_vector(to_unsigned(29, 8)),
			2754 => std_logic_vector(to_unsigned(242, 8)),
			2755 => std_logic_vector(to_unsigned(124, 8)),
			2756 => std_logic_vector(to_unsigned(251, 8)),
			2757 => std_logic_vector(to_unsigned(80, 8)),
			2758 => std_logic_vector(to_unsigned(8, 8)),
			2759 => std_logic_vector(to_unsigned(106, 8)),
			2760 => std_logic_vector(to_unsigned(129, 8)),
			2761 => std_logic_vector(to_unsigned(37, 8)),
			2762 => std_logic_vector(to_unsigned(21, 8)),
			2763 => std_logic_vector(to_unsigned(114, 8)),
			2764 => std_logic_vector(to_unsigned(253, 8)),
			2765 => std_logic_vector(to_unsigned(50, 8)),
			2766 => std_logic_vector(to_unsigned(114, 8)),
			2767 => std_logic_vector(to_unsigned(122, 8)),
			2768 => std_logic_vector(to_unsigned(129, 8)),
			2769 => std_logic_vector(to_unsigned(213, 8)),
			2770 => std_logic_vector(to_unsigned(153, 8)),
			2771 => std_logic_vector(to_unsigned(64, 8)),
			2772 => std_logic_vector(to_unsigned(192, 8)),
			2773 => std_logic_vector(to_unsigned(149, 8)),
			2774 => std_logic_vector(to_unsigned(78, 8)),
			2775 => std_logic_vector(to_unsigned(84, 8)),
			2776 => std_logic_vector(to_unsigned(62, 8)),
			2777 => std_logic_vector(to_unsigned(96, 8)),
			2778 => std_logic_vector(to_unsigned(221, 8)),
			2779 => std_logic_vector(to_unsigned(68, 8)),
			2780 => std_logic_vector(to_unsigned(17, 8)),
			2781 => std_logic_vector(to_unsigned(252, 8)),
			2782 => std_logic_vector(to_unsigned(149, 8)),
			2783 => std_logic_vector(to_unsigned(45, 8)),
			2784 => std_logic_vector(to_unsigned(153, 8)),
			2785 => std_logic_vector(to_unsigned(240, 8)),
			2786 => std_logic_vector(to_unsigned(80, 8)),
			2787 => std_logic_vector(to_unsigned(144, 8)),
			2788 => std_logic_vector(to_unsigned(128, 8)),
			2789 => std_logic_vector(to_unsigned(22, 8)),
			2790 => std_logic_vector(to_unsigned(168, 8)),
			2791 => std_logic_vector(to_unsigned(231, 8)),
			2792 => std_logic_vector(to_unsigned(103, 8)),
			2793 => std_logic_vector(to_unsigned(164, 8)),
			2794 => std_logic_vector(to_unsigned(174, 8)),
			2795 => std_logic_vector(to_unsigned(3, 8)),
			2796 => std_logic_vector(to_unsigned(143, 8)),
			2797 => std_logic_vector(to_unsigned(91, 8)),
			2798 => std_logic_vector(to_unsigned(4, 8)),
			2799 => std_logic_vector(to_unsigned(191, 8)),
			2800 => std_logic_vector(to_unsigned(92, 8)),
			2801 => std_logic_vector(to_unsigned(91, 8)),
			2802 => std_logic_vector(to_unsigned(129, 8)),
			2803 => std_logic_vector(to_unsigned(248, 8)),
			2804 => std_logic_vector(to_unsigned(50, 8)),
			2805 => std_logic_vector(to_unsigned(81, 8)),
			2806 => std_logic_vector(to_unsigned(88, 8)),
			2807 => std_logic_vector(to_unsigned(79, 8)),
			2808 => std_logic_vector(to_unsigned(164, 8)),
			2809 => std_logic_vector(to_unsigned(208, 8)),
			2810 => std_logic_vector(to_unsigned(173, 8)),
			2811 => std_logic_vector(to_unsigned(227, 8)),
			2812 => std_logic_vector(to_unsigned(119, 8)),
			2813 => std_logic_vector(to_unsigned(249, 8)),
			2814 => std_logic_vector(to_unsigned(136, 8)),
			2815 => std_logic_vector(to_unsigned(132, 8)),
			2816 => std_logic_vector(to_unsigned(200, 8)),
			2817 => std_logic_vector(to_unsigned(129, 8)),
			2818 => std_logic_vector(to_unsigned(148, 8)),
			2819 => std_logic_vector(to_unsigned(85, 8)),
			2820 => std_logic_vector(to_unsigned(81, 8)),
			2821 => std_logic_vector(to_unsigned(150, 8)),
			2822 => std_logic_vector(to_unsigned(187, 8)),
			2823 => std_logic_vector(to_unsigned(77, 8)),
			2824 => std_logic_vector(to_unsigned(12, 8)),
			2825 => std_logic_vector(to_unsigned(211, 8)),
			2826 => std_logic_vector(to_unsigned(112, 8)),
			2827 => std_logic_vector(to_unsigned(168, 8)),
			2828 => std_logic_vector(to_unsigned(119, 8)),
			2829 => std_logic_vector(to_unsigned(122, 8)),
			2830 => std_logic_vector(to_unsigned(58, 8)),
			2831 => std_logic_vector(to_unsigned(224, 8)),
			2832 => std_logic_vector(to_unsigned(128, 8)),
			2833 => std_logic_vector(to_unsigned(142, 8)),
			2834 => std_logic_vector(to_unsigned(232, 8)),
			2835 => std_logic_vector(to_unsigned(210, 8)),
			2836 => std_logic_vector(to_unsigned(172, 8)),
			2837 => std_logic_vector(to_unsigned(189, 8)),
			2838 => std_logic_vector(to_unsigned(158, 8)),
			2839 => std_logic_vector(to_unsigned(134, 8)),
			2840 => std_logic_vector(to_unsigned(30, 8)),
			2841 => std_logic_vector(to_unsigned(135, 8)),
			2842 => std_logic_vector(to_unsigned(214, 8)),
			2843 => std_logic_vector(to_unsigned(191, 8)),
			2844 => std_logic_vector(to_unsigned(126, 8)),
			2845 => std_logic_vector(to_unsigned(16, 8)),
			2846 => std_logic_vector(to_unsigned(125, 8)),
			2847 => std_logic_vector(to_unsigned(156, 8)),
			2848 => std_logic_vector(to_unsigned(90, 8)),
			2849 => std_logic_vector(to_unsigned(149, 8)),
			2850 => std_logic_vector(to_unsigned(175, 8)),
			2851 => std_logic_vector(to_unsigned(151, 8)),
			2852 => std_logic_vector(to_unsigned(255, 8)),
			2853 => std_logic_vector(to_unsigned(119, 8)),
			2854 => std_logic_vector(to_unsigned(247, 8)),
			2855 => std_logic_vector(to_unsigned(172, 8)),
			2856 => std_logic_vector(to_unsigned(178, 8)),
			2857 => std_logic_vector(to_unsigned(62, 8)),
			2858 => std_logic_vector(to_unsigned(236, 8)),
			2859 => std_logic_vector(to_unsigned(74, 8)),
			2860 => std_logic_vector(to_unsigned(184, 8)),
			2861 => std_logic_vector(to_unsigned(45, 8)),
			2862 => std_logic_vector(to_unsigned(126, 8)),
			2863 => std_logic_vector(to_unsigned(238, 8)),
			2864 => std_logic_vector(to_unsigned(82, 8)),
			2865 => std_logic_vector(to_unsigned(221, 8)),
			2866 => std_logic_vector(to_unsigned(174, 8)),
			2867 => std_logic_vector(to_unsigned(243, 8)),
			2868 => std_logic_vector(to_unsigned(167, 8)),
			2869 => std_logic_vector(to_unsigned(230, 8)),
			2870 => std_logic_vector(to_unsigned(167, 8)),
			2871 => std_logic_vector(to_unsigned(21, 8)),
			2872 => std_logic_vector(to_unsigned(240, 8)),
			2873 => std_logic_vector(to_unsigned(115, 8)),
			2874 => std_logic_vector(to_unsigned(165, 8)),
			2875 => std_logic_vector(to_unsigned(48, 8)),
			2876 => std_logic_vector(to_unsigned(188, 8)),
			2877 => std_logic_vector(to_unsigned(193, 8)),
			2878 => std_logic_vector(to_unsigned(216, 8)),
			2879 => std_logic_vector(to_unsigned(91, 8)),
			2880 => std_logic_vector(to_unsigned(201, 8)),
			2881 => std_logic_vector(to_unsigned(154, 8)),
			2882 => std_logic_vector(to_unsigned(72, 8)),
			2883 => std_logic_vector(to_unsigned(64, 8)),
			2884 => std_logic_vector(to_unsigned(78, 8)),
			2885 => std_logic_vector(to_unsigned(1, 8)),
			2886 => std_logic_vector(to_unsigned(19, 8)),
			2887 => std_logic_vector(to_unsigned(255, 8)),
			2888 => std_logic_vector(to_unsigned(191, 8)),
			2889 => std_logic_vector(to_unsigned(253, 8)),
			2890 => std_logic_vector(to_unsigned(62, 8)),
			2891 => std_logic_vector(to_unsigned(193, 8)),
			2892 => std_logic_vector(to_unsigned(89, 8)),
			2893 => std_logic_vector(to_unsigned(109, 8)),
			2894 => std_logic_vector(to_unsigned(151, 8)),
			2895 => std_logic_vector(to_unsigned(90, 8)),
			2896 => std_logic_vector(to_unsigned(135, 8)),
			2897 => std_logic_vector(to_unsigned(42, 8)),
			2898 => std_logic_vector(to_unsigned(237, 8)),
			2899 => std_logic_vector(to_unsigned(140, 8)),
			2900 => std_logic_vector(to_unsigned(252, 8)),
			2901 => std_logic_vector(to_unsigned(92, 8)),
			2902 => std_logic_vector(to_unsigned(205, 8)),
			2903 => std_logic_vector(to_unsigned(19, 8)),
			2904 => std_logic_vector(to_unsigned(217, 8)),
			2905 => std_logic_vector(to_unsigned(199, 8)),
			2906 => std_logic_vector(to_unsigned(129, 8)),
			2907 => std_logic_vector(to_unsigned(104, 8)),
			2908 => std_logic_vector(to_unsigned(195, 8)),
			2909 => std_logic_vector(to_unsigned(27, 8)),
			2910 => std_logic_vector(to_unsigned(67, 8)),
			2911 => std_logic_vector(to_unsigned(147, 8)),
			2912 => std_logic_vector(to_unsigned(60, 8)),
			2913 => std_logic_vector(to_unsigned(91, 8)),
			2914 => std_logic_vector(to_unsigned(191, 8)),
			2915 => std_logic_vector(to_unsigned(14, 8)),
			2916 => std_logic_vector(to_unsigned(14, 8)),
			2917 => std_logic_vector(to_unsigned(178, 8)),
			2918 => std_logic_vector(to_unsigned(111, 8)),
			2919 => std_logic_vector(to_unsigned(25, 8)),
			2920 => std_logic_vector(to_unsigned(3, 8)),
			2921 => std_logic_vector(to_unsigned(105, 8)),
			2922 => std_logic_vector(to_unsigned(166, 8)),
			2923 => std_logic_vector(to_unsigned(9, 8)),
			2924 => std_logic_vector(to_unsigned(75, 8)),
			2925 => std_logic_vector(to_unsigned(119, 8)),
			2926 => std_logic_vector(to_unsigned(40, 8)),
			2927 => std_logic_vector(to_unsigned(195, 8)),
			2928 => std_logic_vector(to_unsigned(70, 8)),
			2929 => std_logic_vector(to_unsigned(105, 8)),
			2930 => std_logic_vector(to_unsigned(194, 8)),
			2931 => std_logic_vector(to_unsigned(30, 8)),
			2932 => std_logic_vector(to_unsigned(216, 8)),
			2933 => std_logic_vector(to_unsigned(201, 8)),
			2934 => std_logic_vector(to_unsigned(160, 8)),
			2935 => std_logic_vector(to_unsigned(161, 8)),
			2936 => std_logic_vector(to_unsigned(187, 8)),
			2937 => std_logic_vector(to_unsigned(146, 8)),
			2938 => std_logic_vector(to_unsigned(145, 8)),
			2939 => std_logic_vector(to_unsigned(72, 8)),
			2940 => std_logic_vector(to_unsigned(47, 8)),
			2941 => std_logic_vector(to_unsigned(133, 8)),
			2942 => std_logic_vector(to_unsigned(211, 8)),
			2943 => std_logic_vector(to_unsigned(249, 8)),
			2944 => std_logic_vector(to_unsigned(158, 8)),
			2945 => std_logic_vector(to_unsigned(81, 8)),
			2946 => std_logic_vector(to_unsigned(237, 8)),
			2947 => std_logic_vector(to_unsigned(154, 8)),
			2948 => std_logic_vector(to_unsigned(241, 8)),
			2949 => std_logic_vector(to_unsigned(246, 8)),
			2950 => std_logic_vector(to_unsigned(128, 8)),
			2951 => std_logic_vector(to_unsigned(180, 8)),
			2952 => std_logic_vector(to_unsigned(115, 8)),
			2953 => std_logic_vector(to_unsigned(151, 8)),
			2954 => std_logic_vector(to_unsigned(225, 8)),
			2955 => std_logic_vector(to_unsigned(124, 8)),
			2956 => std_logic_vector(to_unsigned(10, 8)),
			2957 => std_logic_vector(to_unsigned(226, 8)),
			2958 => std_logic_vector(to_unsigned(136, 8)),
			2959 => std_logic_vector(to_unsigned(84, 8)),
			2960 => std_logic_vector(to_unsigned(238, 8)),
			2961 => std_logic_vector(to_unsigned(177, 8)),
			2962 => std_logic_vector(to_unsigned(127, 8)),
			2963 => std_logic_vector(to_unsigned(104, 8)),
			2964 => std_logic_vector(to_unsigned(248, 8)),
			2965 => std_logic_vector(to_unsigned(163, 8)),
			2966 => std_logic_vector(to_unsigned(78, 8)),
			2967 => std_logic_vector(to_unsigned(16, 8)),
			2968 => std_logic_vector(to_unsigned(5, 8)),
			2969 => std_logic_vector(to_unsigned(17, 8)),
			2970 => std_logic_vector(to_unsigned(19, 8)),
			2971 => std_logic_vector(to_unsigned(187, 8)),
			2972 => std_logic_vector(to_unsigned(58, 8)),
			2973 => std_logic_vector(to_unsigned(83, 8)),
			2974 => std_logic_vector(to_unsigned(26, 8)),
			2975 => std_logic_vector(to_unsigned(203, 8)),
			2976 => std_logic_vector(to_unsigned(42, 8)),
			2977 => std_logic_vector(to_unsigned(229, 8)),
			2978 => std_logic_vector(to_unsigned(91, 8)),
			2979 => std_logic_vector(to_unsigned(163, 8)),
			2980 => std_logic_vector(to_unsigned(249, 8)),
			2981 => std_logic_vector(to_unsigned(173, 8)),
			2982 => std_logic_vector(to_unsigned(128, 8)),
			2983 => std_logic_vector(to_unsigned(73, 8)),
			2984 => std_logic_vector(to_unsigned(155, 8)),
			2985 => std_logic_vector(to_unsigned(248, 8)),
			2986 => std_logic_vector(to_unsigned(120, 8)),
			2987 => std_logic_vector(to_unsigned(119, 8)),
			2988 => std_logic_vector(to_unsigned(220, 8)),
			2989 => std_logic_vector(to_unsigned(239, 8)),
			2990 => std_logic_vector(to_unsigned(184, 8)),
			2991 => std_logic_vector(to_unsigned(121, 8)),
			2992 => std_logic_vector(to_unsigned(210, 8)),
			2993 => std_logic_vector(to_unsigned(187, 8)),
			2994 => std_logic_vector(to_unsigned(225, 8)),
			2995 => std_logic_vector(to_unsigned(76, 8)),
			2996 => std_logic_vector(to_unsigned(128, 8)),
			2997 => std_logic_vector(to_unsigned(15, 8)),
			2998 => std_logic_vector(to_unsigned(0, 8)),
			2999 => std_logic_vector(to_unsigned(25, 8)),
			3000 => std_logic_vector(to_unsigned(192, 8)),
			3001 => std_logic_vector(to_unsigned(16, 8)),
			3002 => std_logic_vector(to_unsigned(18, 8)),
			3003 => std_logic_vector(to_unsigned(255, 8)),
			3004 => std_logic_vector(to_unsigned(220, 8)),
			3005 => std_logic_vector(to_unsigned(5, 8)),
			3006 => std_logic_vector(to_unsigned(78, 8)),
			3007 => std_logic_vector(to_unsigned(232, 8)),
			3008 => std_logic_vector(to_unsigned(224, 8)),
			3009 => std_logic_vector(to_unsigned(124, 8)),
			3010 => std_logic_vector(to_unsigned(7, 8)),
			3011 => std_logic_vector(to_unsigned(22, 8)),
			3012 => std_logic_vector(to_unsigned(34, 8)),
			3013 => std_logic_vector(to_unsigned(241, 8)),
			3014 => std_logic_vector(to_unsigned(244, 8)),
			3015 => std_logic_vector(to_unsigned(75, 8)),
			3016 => std_logic_vector(to_unsigned(218, 8)),
			3017 => std_logic_vector(to_unsigned(121, 8)),
			3018 => std_logic_vector(to_unsigned(232, 8)),
			3019 => std_logic_vector(to_unsigned(13, 8)),
			3020 => std_logic_vector(to_unsigned(0, 8)),
			3021 => std_logic_vector(to_unsigned(98, 8)),
			3022 => std_logic_vector(to_unsigned(179, 8)),
			3023 => std_logic_vector(to_unsigned(79, 8)),
			3024 => std_logic_vector(to_unsigned(173, 8)),
			3025 => std_logic_vector(to_unsigned(59, 8)),
			3026 => std_logic_vector(to_unsigned(55, 8)),
			3027 => std_logic_vector(to_unsigned(40, 8)),
			3028 => std_logic_vector(to_unsigned(89, 8)),
			3029 => std_logic_vector(to_unsigned(87, 8)),
			3030 => std_logic_vector(to_unsigned(201, 8)),
			3031 => std_logic_vector(to_unsigned(75, 8)),
			3032 => std_logic_vector(to_unsigned(24, 8)),
			3033 => std_logic_vector(to_unsigned(161, 8)),
			3034 => std_logic_vector(to_unsigned(211, 8)),
			3035 => std_logic_vector(to_unsigned(78, 8)),
			3036 => std_logic_vector(to_unsigned(176, 8)),
			3037 => std_logic_vector(to_unsigned(113, 8)),
			3038 => std_logic_vector(to_unsigned(207, 8)),
			3039 => std_logic_vector(to_unsigned(231, 8)),
			3040 => std_logic_vector(to_unsigned(78, 8)),
			3041 => std_logic_vector(to_unsigned(186, 8)),
			3042 => std_logic_vector(to_unsigned(95, 8)),
			3043 => std_logic_vector(to_unsigned(6, 8)),
			3044 => std_logic_vector(to_unsigned(244, 8)),
			3045 => std_logic_vector(to_unsigned(46, 8)),
			3046 => std_logic_vector(to_unsigned(51, 8)),
			3047 => std_logic_vector(to_unsigned(216, 8)),
			3048 => std_logic_vector(to_unsigned(203, 8)),
			3049 => std_logic_vector(to_unsigned(2, 8)),
			3050 => std_logic_vector(to_unsigned(10, 8)),
			3051 => std_logic_vector(to_unsigned(216, 8)),
			3052 => std_logic_vector(to_unsigned(117, 8)),
			3053 => std_logic_vector(to_unsigned(29, 8)),
			3054 => std_logic_vector(to_unsigned(45, 8)),
			3055 => std_logic_vector(to_unsigned(48, 8)),
			3056 => std_logic_vector(to_unsigned(97, 8)),
			3057 => std_logic_vector(to_unsigned(124, 8)),
			3058 => std_logic_vector(to_unsigned(22, 8)),
			3059 => std_logic_vector(to_unsigned(146, 8)),
			3060 => std_logic_vector(to_unsigned(138, 8)),
			3061 => std_logic_vector(to_unsigned(140, 8)),
			3062 => std_logic_vector(to_unsigned(204, 8)),
			3063 => std_logic_vector(to_unsigned(94, 8)),
			3064 => std_logic_vector(to_unsigned(231, 8)),
			3065 => std_logic_vector(to_unsigned(119, 8)),
			3066 => std_logic_vector(to_unsigned(111, 8)),
			3067 => std_logic_vector(to_unsigned(137, 8)),
			3068 => std_logic_vector(to_unsigned(162, 8)),
			3069 => std_logic_vector(to_unsigned(64, 8)),
			3070 => std_logic_vector(to_unsigned(22, 8)),
			3071 => std_logic_vector(to_unsigned(225, 8)),
			3072 => std_logic_vector(to_unsigned(103, 8)),
			3073 => std_logic_vector(to_unsigned(226, 8)),
			3074 => std_logic_vector(to_unsigned(113, 8)),
			3075 => std_logic_vector(to_unsigned(143, 8)),
			3076 => std_logic_vector(to_unsigned(98, 8)),
			3077 => std_logic_vector(to_unsigned(225, 8)),
			3078 => std_logic_vector(to_unsigned(133, 8)),
			3079 => std_logic_vector(to_unsigned(207, 8)),
			3080 => std_logic_vector(to_unsigned(224, 8)),
			3081 => std_logic_vector(to_unsigned(112, 8)),
			3082 => std_logic_vector(to_unsigned(254, 8)),
			3083 => std_logic_vector(to_unsigned(49, 8)),
			3084 => std_logic_vector(to_unsigned(54, 8)),
			3085 => std_logic_vector(to_unsigned(157, 8)),
			3086 => std_logic_vector(to_unsigned(179, 8)),
			3087 => std_logic_vector(to_unsigned(217, 8)),
			3088 => std_logic_vector(to_unsigned(235, 8)),
			3089 => std_logic_vector(to_unsigned(214, 8)),
			3090 => std_logic_vector(to_unsigned(70, 8)),
			3091 => std_logic_vector(to_unsigned(36, 8)),
			3092 => std_logic_vector(to_unsigned(81, 8)),
			3093 => std_logic_vector(to_unsigned(213, 8)),
			3094 => std_logic_vector(to_unsigned(174, 8)),
			3095 => std_logic_vector(to_unsigned(209, 8)),
			3096 => std_logic_vector(to_unsigned(202, 8)),
			3097 => std_logic_vector(to_unsigned(112, 8)),
			3098 => std_logic_vector(to_unsigned(122, 8)),
			3099 => std_logic_vector(to_unsigned(159, 8)),
			3100 => std_logic_vector(to_unsigned(243, 8)),
			3101 => std_logic_vector(to_unsigned(21, 8)),
			3102 => std_logic_vector(to_unsigned(19, 8)),
			3103 => std_logic_vector(to_unsigned(151, 8)),
			3104 => std_logic_vector(to_unsigned(48, 8)),
			3105 => std_logic_vector(to_unsigned(239, 8)),
			3106 => std_logic_vector(to_unsigned(255, 8)),
			3107 => std_logic_vector(to_unsigned(116, 8)),
			3108 => std_logic_vector(to_unsigned(107, 8)),
			3109 => std_logic_vector(to_unsigned(145, 8)),
			3110 => std_logic_vector(to_unsigned(62, 8)),
			3111 => std_logic_vector(to_unsigned(109, 8)),
			3112 => std_logic_vector(to_unsigned(28, 8)),
			3113 => std_logic_vector(to_unsigned(193, 8)),
			3114 => std_logic_vector(to_unsigned(94, 8)),
			3115 => std_logic_vector(to_unsigned(169, 8)),
			3116 => std_logic_vector(to_unsigned(13, 8)),
			3117 => std_logic_vector(to_unsigned(136, 8)),
			3118 => std_logic_vector(to_unsigned(36, 8)),
			3119 => std_logic_vector(to_unsigned(168, 8)),
			3120 => std_logic_vector(to_unsigned(111, 8)),
			3121 => std_logic_vector(to_unsigned(121, 8)),
			3122 => std_logic_vector(to_unsigned(238, 8)),
			3123 => std_logic_vector(to_unsigned(142, 8)),
			3124 => std_logic_vector(to_unsigned(231, 8)),
			3125 => std_logic_vector(to_unsigned(206, 8)),
			3126 => std_logic_vector(to_unsigned(209, 8)),
			3127 => std_logic_vector(to_unsigned(62, 8)),
			3128 => std_logic_vector(to_unsigned(192, 8)),
			3129 => std_logic_vector(to_unsigned(15, 8)),
			3130 => std_logic_vector(to_unsigned(178, 8)),
			3131 => std_logic_vector(to_unsigned(51, 8)),
			3132 => std_logic_vector(to_unsigned(17, 8)),
			3133 => std_logic_vector(to_unsigned(34, 8)),
			3134 => std_logic_vector(to_unsigned(156, 8)),
			3135 => std_logic_vector(to_unsigned(128, 8)),
			3136 => std_logic_vector(to_unsigned(201, 8)),
			3137 => std_logic_vector(to_unsigned(217, 8)),
			3138 => std_logic_vector(to_unsigned(12, 8)),
			3139 => std_logic_vector(to_unsigned(20, 8)),
			3140 => std_logic_vector(to_unsigned(146, 8)),
			3141 => std_logic_vector(to_unsigned(212, 8)),
			3142 => std_logic_vector(to_unsigned(151, 8)),
			3143 => std_logic_vector(to_unsigned(112, 8)),
			3144 => std_logic_vector(to_unsigned(127, 8)),
			3145 => std_logic_vector(to_unsigned(223, 8)),
			3146 => std_logic_vector(to_unsigned(112, 8)),
			3147 => std_logic_vector(to_unsigned(147, 8)),
			3148 => std_logic_vector(to_unsigned(140, 8)),
			3149 => std_logic_vector(to_unsigned(217, 8)),
			3150 => std_logic_vector(to_unsigned(167, 8)),
			3151 => std_logic_vector(to_unsigned(142, 8)),
			3152 => std_logic_vector(to_unsigned(161, 8)),
			3153 => std_logic_vector(to_unsigned(84, 8)),
			3154 => std_logic_vector(to_unsigned(199, 8)),
			3155 => std_logic_vector(to_unsigned(173, 8)),
			3156 => std_logic_vector(to_unsigned(31, 8)),
			3157 => std_logic_vector(to_unsigned(121, 8)),
			3158 => std_logic_vector(to_unsigned(126, 8)),
			3159 => std_logic_vector(to_unsigned(106, 8)),
			3160 => std_logic_vector(to_unsigned(57, 8)),
			3161 => std_logic_vector(to_unsigned(172, 8)),
			3162 => std_logic_vector(to_unsigned(185, 8)),
			3163 => std_logic_vector(to_unsigned(124, 8)),
			3164 => std_logic_vector(to_unsigned(62, 8)),
			3165 => std_logic_vector(to_unsigned(237, 8)),
			3166 => std_logic_vector(to_unsigned(87, 8)),
			3167 => std_logic_vector(to_unsigned(187, 8)),
			3168 => std_logic_vector(to_unsigned(173, 8)),
			3169 => std_logic_vector(to_unsigned(238, 8)),
			3170 => std_logic_vector(to_unsigned(214, 8)),
			3171 => std_logic_vector(to_unsigned(149, 8)),
			3172 => std_logic_vector(to_unsigned(54, 8)),
			3173 => std_logic_vector(to_unsigned(219, 8)),
			3174 => std_logic_vector(to_unsigned(23, 8)),
			3175 => std_logic_vector(to_unsigned(244, 8)),
			3176 => std_logic_vector(to_unsigned(181, 8)),
			3177 => std_logic_vector(to_unsigned(147, 8)),
			3178 => std_logic_vector(to_unsigned(41, 8)),
			3179 => std_logic_vector(to_unsigned(204, 8)),
			3180 => std_logic_vector(to_unsigned(133, 8)),
			3181 => std_logic_vector(to_unsigned(91, 8)),
			3182 => std_logic_vector(to_unsigned(29, 8)),
			3183 => std_logic_vector(to_unsigned(165, 8)),
			3184 => std_logic_vector(to_unsigned(107, 8)),
			3185 => std_logic_vector(to_unsigned(141, 8)),
			3186 => std_logic_vector(to_unsigned(145, 8)),
			3187 => std_logic_vector(to_unsigned(117, 8)),
			3188 => std_logic_vector(to_unsigned(32, 8)),
			3189 => std_logic_vector(to_unsigned(89, 8)),
			3190 => std_logic_vector(to_unsigned(191, 8)),
			3191 => std_logic_vector(to_unsigned(190, 8)),
			3192 => std_logic_vector(to_unsigned(83, 8)),
			3193 => std_logic_vector(to_unsigned(214, 8)),
			3194 => std_logic_vector(to_unsigned(219, 8)),
			3195 => std_logic_vector(to_unsigned(144, 8)),
			3196 => std_logic_vector(to_unsigned(241, 8)),
			3197 => std_logic_vector(to_unsigned(114, 8)),
			3198 => std_logic_vector(to_unsigned(250, 8)),
			3199 => std_logic_vector(to_unsigned(69, 8)),
			3200 => std_logic_vector(to_unsigned(93, 8)),
			3201 => std_logic_vector(to_unsigned(45, 8)),
			3202 => std_logic_vector(to_unsigned(82, 8)),
			3203 => std_logic_vector(to_unsigned(97, 8)),
			3204 => std_logic_vector(to_unsigned(140, 8)),
			3205 => std_logic_vector(to_unsigned(32, 8)),
			3206 => std_logic_vector(to_unsigned(60, 8)),
			3207 => std_logic_vector(to_unsigned(14, 8)),
			3208 => std_logic_vector(to_unsigned(148, 8)),
			3209 => std_logic_vector(to_unsigned(31, 8)),
			3210 => std_logic_vector(to_unsigned(45, 8)),
			3211 => std_logic_vector(to_unsigned(164, 8)),
			3212 => std_logic_vector(to_unsigned(66, 8)),
			3213 => std_logic_vector(to_unsigned(77, 8)),
			3214 => std_logic_vector(to_unsigned(51, 8)),
			3215 => std_logic_vector(to_unsigned(139, 8)),
			3216 => std_logic_vector(to_unsigned(17, 8)),
			3217 => std_logic_vector(to_unsigned(228, 8)),
			3218 => std_logic_vector(to_unsigned(57, 8)),
			3219 => std_logic_vector(to_unsigned(144, 8)),
			3220 => std_logic_vector(to_unsigned(206, 8)),
			3221 => std_logic_vector(to_unsigned(123, 8)),
			3222 => std_logic_vector(to_unsigned(59, 8)),
			3223 => std_logic_vector(to_unsigned(211, 8)),
			3224 => std_logic_vector(to_unsigned(234, 8)),
			3225 => std_logic_vector(to_unsigned(222, 8)),
			3226 => std_logic_vector(to_unsigned(196, 8)),
			3227 => std_logic_vector(to_unsigned(115, 8)),
			3228 => std_logic_vector(to_unsigned(174, 8)),
			3229 => std_logic_vector(to_unsigned(115, 8)),
			3230 => std_logic_vector(to_unsigned(229, 8)),
			3231 => std_logic_vector(to_unsigned(97, 8)),
			3232 => std_logic_vector(to_unsigned(177, 8)),
			3233 => std_logic_vector(to_unsigned(222, 8)),
			3234 => std_logic_vector(to_unsigned(64, 8)),
			3235 => std_logic_vector(to_unsigned(82, 8)),
			3236 => std_logic_vector(to_unsigned(157, 8)),
			3237 => std_logic_vector(to_unsigned(203, 8)),
			3238 => std_logic_vector(to_unsigned(128, 8)),
			3239 => std_logic_vector(to_unsigned(143, 8)),
			3240 => std_logic_vector(to_unsigned(244, 8)),
			3241 => std_logic_vector(to_unsigned(123, 8)),
			3242 => std_logic_vector(to_unsigned(131, 8)),
			3243 => std_logic_vector(to_unsigned(76, 8)),
			3244 => std_logic_vector(to_unsigned(25, 8)),
			3245 => std_logic_vector(to_unsigned(173, 8)),
			3246 => std_logic_vector(to_unsigned(100, 8)),
			3247 => std_logic_vector(to_unsigned(246, 8)),
			3248 => std_logic_vector(to_unsigned(61, 8)),
			3249 => std_logic_vector(to_unsigned(147, 8)),
			3250 => std_logic_vector(to_unsigned(11, 8)),
			3251 => std_logic_vector(to_unsigned(59, 8)),
			3252 => std_logic_vector(to_unsigned(137, 8)),
			3253 => std_logic_vector(to_unsigned(73, 8)),
			3254 => std_logic_vector(to_unsigned(147, 8)),
			3255 => std_logic_vector(to_unsigned(40, 8)),
			3256 => std_logic_vector(to_unsigned(123, 8)),
			3257 => std_logic_vector(to_unsigned(94, 8)),
			3258 => std_logic_vector(to_unsigned(123, 8)),
			3259 => std_logic_vector(to_unsigned(226, 8)),
			3260 => std_logic_vector(to_unsigned(235, 8)),
			3261 => std_logic_vector(to_unsigned(177, 8)),
			3262 => std_logic_vector(to_unsigned(180, 8)),
			3263 => std_logic_vector(to_unsigned(16, 8)),
			3264 => std_logic_vector(to_unsigned(135, 8)),
			3265 => std_logic_vector(to_unsigned(204, 8)),
			3266 => std_logic_vector(to_unsigned(53, 8)),
			3267 => std_logic_vector(to_unsigned(99, 8)),
			3268 => std_logic_vector(to_unsigned(223, 8)),
			3269 => std_logic_vector(to_unsigned(47, 8)),
			3270 => std_logic_vector(to_unsigned(93, 8)),
			3271 => std_logic_vector(to_unsigned(95, 8)),
			3272 => std_logic_vector(to_unsigned(168, 8)),
			3273 => std_logic_vector(to_unsigned(207, 8)),
			3274 => std_logic_vector(to_unsigned(36, 8)),
			3275 => std_logic_vector(to_unsigned(45, 8)),
			3276 => std_logic_vector(to_unsigned(131, 8)),
			3277 => std_logic_vector(to_unsigned(251, 8)),
			3278 => std_logic_vector(to_unsigned(172, 8)),
			3279 => std_logic_vector(to_unsigned(80, 8)),
			3280 => std_logic_vector(to_unsigned(132, 8)),
			3281 => std_logic_vector(to_unsigned(31, 8)),
			3282 => std_logic_vector(to_unsigned(114, 8)),
			3283 => std_logic_vector(to_unsigned(176, 8)),
			3284 => std_logic_vector(to_unsigned(234, 8)),
			3285 => std_logic_vector(to_unsigned(183, 8)),
			3286 => std_logic_vector(to_unsigned(23, 8)),
			3287 => std_logic_vector(to_unsigned(108, 8)),
			3288 => std_logic_vector(to_unsigned(33, 8)),
			3289 => std_logic_vector(to_unsigned(85, 8)),
			3290 => std_logic_vector(to_unsigned(168, 8)),
			3291 => std_logic_vector(to_unsigned(24, 8)),
			3292 => std_logic_vector(to_unsigned(46, 8)),
			3293 => std_logic_vector(to_unsigned(23, 8)),
			3294 => std_logic_vector(to_unsigned(180, 8)),
			3295 => std_logic_vector(to_unsigned(111, 8)),
			3296 => std_logic_vector(to_unsigned(75, 8)),
			3297 => std_logic_vector(to_unsigned(166, 8)),
			3298 => std_logic_vector(to_unsigned(172, 8)),
			3299 => std_logic_vector(to_unsigned(26, 8)),
			3300 => std_logic_vector(to_unsigned(54, 8)),
			3301 => std_logic_vector(to_unsigned(171, 8)),
			3302 => std_logic_vector(to_unsigned(66, 8)),
			3303 => std_logic_vector(to_unsigned(179, 8)),
			3304 => std_logic_vector(to_unsigned(98, 8)),
			3305 => std_logic_vector(to_unsigned(199, 8)),
			3306 => std_logic_vector(to_unsigned(155, 8)),
			3307 => std_logic_vector(to_unsigned(88, 8)),
			3308 => std_logic_vector(to_unsigned(91, 8)),
			3309 => std_logic_vector(to_unsigned(134, 8)),
			3310 => std_logic_vector(to_unsigned(49, 8)),
			3311 => std_logic_vector(to_unsigned(49, 8)),
			3312 => std_logic_vector(to_unsigned(54, 8)),
			3313 => std_logic_vector(to_unsigned(146, 8)),
			3314 => std_logic_vector(to_unsigned(19, 8)),
			3315 => std_logic_vector(to_unsigned(181, 8)),
			3316 => std_logic_vector(to_unsigned(201, 8)),
			3317 => std_logic_vector(to_unsigned(121, 8)),
			3318 => std_logic_vector(to_unsigned(109, 8)),
			3319 => std_logic_vector(to_unsigned(109, 8)),
			3320 => std_logic_vector(to_unsigned(32, 8)),
			3321 => std_logic_vector(to_unsigned(12, 8)),
			3322 => std_logic_vector(to_unsigned(80, 8)),
			3323 => std_logic_vector(to_unsigned(176, 8)),
			3324 => std_logic_vector(to_unsigned(208, 8)),
			3325 => std_logic_vector(to_unsigned(139, 8)),
			3326 => std_logic_vector(to_unsigned(199, 8)),
			3327 => std_logic_vector(to_unsigned(194, 8)),
			3328 => std_logic_vector(to_unsigned(244, 8)),
			3329 => std_logic_vector(to_unsigned(23, 8)),
			3330 => std_logic_vector(to_unsigned(93, 8)),
			3331 => std_logic_vector(to_unsigned(138, 8)),
			3332 => std_logic_vector(to_unsigned(208, 8)),
			3333 => std_logic_vector(to_unsigned(126, 8)),
			3334 => std_logic_vector(to_unsigned(200, 8)),
			3335 => std_logic_vector(to_unsigned(8, 8)),
			3336 => std_logic_vector(to_unsigned(236, 8)),
			3337 => std_logic_vector(to_unsigned(97, 8)),
			3338 => std_logic_vector(to_unsigned(74, 8)),
			3339 => std_logic_vector(to_unsigned(12, 8)),
			3340 => std_logic_vector(to_unsigned(84, 8)),
			3341 => std_logic_vector(to_unsigned(119, 8)),
			3342 => std_logic_vector(to_unsigned(18, 8)),
			3343 => std_logic_vector(to_unsigned(210, 8)),
			3344 => std_logic_vector(to_unsigned(42, 8)),
			3345 => std_logic_vector(to_unsigned(50, 8)),
			3346 => std_logic_vector(to_unsigned(29, 8)),
			3347 => std_logic_vector(to_unsigned(234, 8)),
			3348 => std_logic_vector(to_unsigned(57, 8)),
			3349 => std_logic_vector(to_unsigned(105, 8)),
			3350 => std_logic_vector(to_unsigned(164, 8)),
			3351 => std_logic_vector(to_unsigned(76, 8)),
			3352 => std_logic_vector(to_unsigned(172, 8)),
			3353 => std_logic_vector(to_unsigned(30, 8)),
			3354 => std_logic_vector(to_unsigned(108, 8)),
			3355 => std_logic_vector(to_unsigned(163, 8)),
			3356 => std_logic_vector(to_unsigned(8, 8)),
			3357 => std_logic_vector(to_unsigned(113, 8)),
			3358 => std_logic_vector(to_unsigned(218, 8)),
			3359 => std_logic_vector(to_unsigned(179, 8)),
			3360 => std_logic_vector(to_unsigned(214, 8)),
			3361 => std_logic_vector(to_unsigned(232, 8)),
			3362 => std_logic_vector(to_unsigned(36, 8)),
			3363 => std_logic_vector(to_unsigned(27, 8)),
			3364 => std_logic_vector(to_unsigned(129, 8)),
			3365 => std_logic_vector(to_unsigned(244, 8)),
			3366 => std_logic_vector(to_unsigned(90, 8)),
			3367 => std_logic_vector(to_unsigned(20, 8)),
			3368 => std_logic_vector(to_unsigned(51, 8)),
			3369 => std_logic_vector(to_unsigned(79, 8)),
			3370 => std_logic_vector(to_unsigned(63, 8)),
			3371 => std_logic_vector(to_unsigned(234, 8)),
			3372 => std_logic_vector(to_unsigned(67, 8)),
			3373 => std_logic_vector(to_unsigned(137, 8)),
			3374 => std_logic_vector(to_unsigned(57, 8)),
			3375 => std_logic_vector(to_unsigned(133, 8)),
			3376 => std_logic_vector(to_unsigned(8, 8)),
			3377 => std_logic_vector(to_unsigned(86, 8)),
			3378 => std_logic_vector(to_unsigned(254, 8)),
			3379 => std_logic_vector(to_unsigned(181, 8)),
			3380 => std_logic_vector(to_unsigned(126, 8)),
			3381 => std_logic_vector(to_unsigned(173, 8)),
			3382 => std_logic_vector(to_unsigned(45, 8)),
			3383 => std_logic_vector(to_unsigned(35, 8)),
			3384 => std_logic_vector(to_unsigned(198, 8)),
			3385 => std_logic_vector(to_unsigned(152, 8)),
			3386 => std_logic_vector(to_unsigned(173, 8)),
			3387 => std_logic_vector(to_unsigned(83, 8)),
			3388 => std_logic_vector(to_unsigned(10, 8)),
			3389 => std_logic_vector(to_unsigned(132, 8)),
			3390 => std_logic_vector(to_unsigned(164, 8)),
			3391 => std_logic_vector(to_unsigned(127, 8)),
			3392 => std_logic_vector(to_unsigned(54, 8)),
			3393 => std_logic_vector(to_unsigned(237, 8)),
			3394 => std_logic_vector(to_unsigned(248, 8)),
			3395 => std_logic_vector(to_unsigned(115, 8)),
			3396 => std_logic_vector(to_unsigned(102, 8)),
			3397 => std_logic_vector(to_unsigned(86, 8)),
			3398 => std_logic_vector(to_unsigned(232, 8)),
			3399 => std_logic_vector(to_unsigned(46, 8)),
			3400 => std_logic_vector(to_unsigned(148, 8)),
			3401 => std_logic_vector(to_unsigned(78, 8)),
			3402 => std_logic_vector(to_unsigned(79, 8)),
			3403 => std_logic_vector(to_unsigned(126, 8)),
			3404 => std_logic_vector(to_unsigned(97, 8)),
			3405 => std_logic_vector(to_unsigned(143, 8)),
			3406 => std_logic_vector(to_unsigned(133, 8)),
			3407 => std_logic_vector(to_unsigned(11, 8)),
			3408 => std_logic_vector(to_unsigned(156, 8)),
			3409 => std_logic_vector(to_unsigned(187, 8)),
			3410 => std_logic_vector(to_unsigned(184, 8)),
			3411 => std_logic_vector(to_unsigned(97, 8)),
			3412 => std_logic_vector(to_unsigned(151, 8)),
			3413 => std_logic_vector(to_unsigned(237, 8)),
			3414 => std_logic_vector(to_unsigned(49, 8)),
			3415 => std_logic_vector(to_unsigned(42, 8)),
			3416 => std_logic_vector(to_unsigned(21, 8)),
			3417 => std_logic_vector(to_unsigned(177, 8)),
			3418 => std_logic_vector(to_unsigned(55, 8)),
			3419 => std_logic_vector(to_unsigned(111, 8)),
			3420 => std_logic_vector(to_unsigned(2, 8)),
			3421 => std_logic_vector(to_unsigned(246, 8)),
			3422 => std_logic_vector(to_unsigned(101, 8)),
			3423 => std_logic_vector(to_unsigned(131, 8)),
			3424 => std_logic_vector(to_unsigned(14, 8)),
			3425 => std_logic_vector(to_unsigned(159, 8)),
			3426 => std_logic_vector(to_unsigned(210, 8)),
			3427 => std_logic_vector(to_unsigned(174, 8)),
			3428 => std_logic_vector(to_unsigned(204, 8)),
			3429 => std_logic_vector(to_unsigned(109, 8)),
			3430 => std_logic_vector(to_unsigned(242, 8)),
			3431 => std_logic_vector(to_unsigned(114, 8)),
			3432 => std_logic_vector(to_unsigned(219, 8)),
			3433 => std_logic_vector(to_unsigned(29, 8)),
			3434 => std_logic_vector(to_unsigned(84, 8)),
			3435 => std_logic_vector(to_unsigned(113, 8)),
			3436 => std_logic_vector(to_unsigned(85, 8)),
			3437 => std_logic_vector(to_unsigned(177, 8)),
			3438 => std_logic_vector(to_unsigned(163, 8)),
			3439 => std_logic_vector(to_unsigned(188, 8)),
			3440 => std_logic_vector(to_unsigned(249, 8)),
			3441 => std_logic_vector(to_unsigned(10, 8)),
			3442 => std_logic_vector(to_unsigned(68, 8)),
			3443 => std_logic_vector(to_unsigned(2, 8)),
			3444 => std_logic_vector(to_unsigned(235, 8)),
			3445 => std_logic_vector(to_unsigned(97, 8)),
			3446 => std_logic_vector(to_unsigned(226, 8)),
			3447 => std_logic_vector(to_unsigned(87, 8)),
			3448 => std_logic_vector(to_unsigned(52, 8)),
			3449 => std_logic_vector(to_unsigned(44, 8)),
			3450 => std_logic_vector(to_unsigned(180, 8)),
			3451 => std_logic_vector(to_unsigned(40, 8)),
			3452 => std_logic_vector(to_unsigned(96, 8)),
			3453 => std_logic_vector(to_unsigned(99, 8)),
			3454 => std_logic_vector(to_unsigned(63, 8)),
			3455 => std_logic_vector(to_unsigned(204, 8)),
			3456 => std_logic_vector(to_unsigned(85, 8)),
			3457 => std_logic_vector(to_unsigned(93, 8)),
			3458 => std_logic_vector(to_unsigned(67, 8)),
			3459 => std_logic_vector(to_unsigned(252, 8)),
			3460 => std_logic_vector(to_unsigned(241, 8)),
			3461 => std_logic_vector(to_unsigned(6, 8)),
			3462 => std_logic_vector(to_unsigned(232, 8)),
			3463 => std_logic_vector(to_unsigned(222, 8)),
			3464 => std_logic_vector(to_unsigned(191, 8)),
			3465 => std_logic_vector(to_unsigned(146, 8)),
			3466 => std_logic_vector(to_unsigned(220, 8)),
			3467 => std_logic_vector(to_unsigned(150, 8)),
			3468 => std_logic_vector(to_unsigned(192, 8)),
			3469 => std_logic_vector(to_unsigned(88, 8)),
			3470 => std_logic_vector(to_unsigned(235, 8)),
			3471 => std_logic_vector(to_unsigned(145, 8)),
			3472 => std_logic_vector(to_unsigned(198, 8)),
			3473 => std_logic_vector(to_unsigned(90, 8)),
			3474 => std_logic_vector(to_unsigned(154, 8)),
			3475 => std_logic_vector(to_unsigned(38, 8)),
			3476 => std_logic_vector(to_unsigned(177, 8)),
			3477 => std_logic_vector(to_unsigned(236, 8)),
			3478 => std_logic_vector(to_unsigned(197, 8)),
			3479 => std_logic_vector(to_unsigned(202, 8)),
			3480 => std_logic_vector(to_unsigned(193, 8)),
			3481 => std_logic_vector(to_unsigned(220, 8)),
			3482 => std_logic_vector(to_unsigned(173, 8)),
			3483 => std_logic_vector(to_unsigned(241, 8)),
			3484 => std_logic_vector(to_unsigned(230, 8)),
			3485 => std_logic_vector(to_unsigned(250, 8)),
			3486 => std_logic_vector(to_unsigned(185, 8)),
			3487 => std_logic_vector(to_unsigned(32, 8)),
			3488 => std_logic_vector(to_unsigned(152, 8)),
			3489 => std_logic_vector(to_unsigned(1, 8)),
			3490 => std_logic_vector(to_unsigned(218, 8)),
			3491 => std_logic_vector(to_unsigned(235, 8)),
			3492 => std_logic_vector(to_unsigned(189, 8)),
			3493 => std_logic_vector(to_unsigned(147, 8)),
			3494 => std_logic_vector(to_unsigned(207, 8)),
			3495 => std_logic_vector(to_unsigned(49, 8)),
			3496 => std_logic_vector(to_unsigned(3, 8)),
			3497 => std_logic_vector(to_unsigned(136, 8)),
			3498 => std_logic_vector(to_unsigned(245, 8)),
			3499 => std_logic_vector(to_unsigned(110, 8)),
			3500 => std_logic_vector(to_unsigned(151, 8)),
			3501 => std_logic_vector(to_unsigned(29, 8)),
			3502 => std_logic_vector(to_unsigned(67, 8)),
			3503 => std_logic_vector(to_unsigned(84, 8)),
			3504 => std_logic_vector(to_unsigned(69, 8)),
			3505 => std_logic_vector(to_unsigned(99, 8)),
			3506 => std_logic_vector(to_unsigned(171, 8)),
			3507 => std_logic_vector(to_unsigned(164, 8)),
			3508 => std_logic_vector(to_unsigned(109, 8)),
			3509 => std_logic_vector(to_unsigned(4, 8)),
			3510 => std_logic_vector(to_unsigned(177, 8)),
			3511 => std_logic_vector(to_unsigned(81, 8)),
			3512 => std_logic_vector(to_unsigned(176, 8)),
			3513 => std_logic_vector(to_unsigned(196, 8)),
			3514 => std_logic_vector(to_unsigned(109, 8)),
			3515 => std_logic_vector(to_unsigned(122, 8)),
			3516 => std_logic_vector(to_unsigned(142, 8)),
			3517 => std_logic_vector(to_unsigned(228, 8)),
			3518 => std_logic_vector(to_unsigned(58, 8)),
			3519 => std_logic_vector(to_unsigned(61, 8)),
			3520 => std_logic_vector(to_unsigned(176, 8)),
			3521 => std_logic_vector(to_unsigned(222, 8)),
			3522 => std_logic_vector(to_unsigned(192, 8)),
			3523 => std_logic_vector(to_unsigned(38, 8)),
			3524 => std_logic_vector(to_unsigned(106, 8)),
			3525 => std_logic_vector(to_unsigned(6, 8)),
			3526 => std_logic_vector(to_unsigned(106, 8)),
			3527 => std_logic_vector(to_unsigned(190, 8)),
			3528 => std_logic_vector(to_unsigned(105, 8)),
			3529 => std_logic_vector(to_unsigned(24, 8)),
			3530 => std_logic_vector(to_unsigned(238, 8)),
			3531 => std_logic_vector(to_unsigned(178, 8)),
			3532 => std_logic_vector(to_unsigned(29, 8)),
			3533 => std_logic_vector(to_unsigned(251, 8)),
			3534 => std_logic_vector(to_unsigned(79, 8)),
			3535 => std_logic_vector(to_unsigned(170, 8)),
			3536 => std_logic_vector(to_unsigned(169, 8)),
			3537 => std_logic_vector(to_unsigned(183, 8)),
			3538 => std_logic_vector(to_unsigned(137, 8)),
			3539 => std_logic_vector(to_unsigned(64, 8)),
			3540 => std_logic_vector(to_unsigned(94, 8)),
			3541 => std_logic_vector(to_unsigned(114, 8)),
			3542 => std_logic_vector(to_unsigned(99, 8)),
			3543 => std_logic_vector(to_unsigned(226, 8)),
			3544 => std_logic_vector(to_unsigned(217, 8)),
			3545 => std_logic_vector(to_unsigned(227, 8)),
			3546 => std_logic_vector(to_unsigned(89, 8)),
			3547 => std_logic_vector(to_unsigned(191, 8)),
			3548 => std_logic_vector(to_unsigned(93, 8)),
			3549 => std_logic_vector(to_unsigned(136, 8)),
			3550 => std_logic_vector(to_unsigned(68, 8)),
			3551 => std_logic_vector(to_unsigned(243, 8)),
			3552 => std_logic_vector(to_unsigned(54, 8)),
			3553 => std_logic_vector(to_unsigned(215, 8)),
			3554 => std_logic_vector(to_unsigned(207, 8)),
			3555 => std_logic_vector(to_unsigned(134, 8)),
			3556 => std_logic_vector(to_unsigned(47, 8)),
			3557 => std_logic_vector(to_unsigned(242, 8)),
			3558 => std_logic_vector(to_unsigned(11, 8)),
			3559 => std_logic_vector(to_unsigned(57, 8)),
			3560 => std_logic_vector(to_unsigned(235, 8)),
			3561 => std_logic_vector(to_unsigned(12, 8)),
			3562 => std_logic_vector(to_unsigned(45, 8)),
			3563 => std_logic_vector(to_unsigned(179, 8)),
			3564 => std_logic_vector(to_unsigned(214, 8)),
			3565 => std_logic_vector(to_unsigned(86, 8)),
			3566 => std_logic_vector(to_unsigned(50, 8)),
			3567 => std_logic_vector(to_unsigned(227, 8)),
			3568 => std_logic_vector(to_unsigned(155, 8)),
			3569 => std_logic_vector(to_unsigned(29, 8)),
			3570 => std_logic_vector(to_unsigned(122, 8)),
			3571 => std_logic_vector(to_unsigned(160, 8)),
			3572 => std_logic_vector(to_unsigned(154, 8)),
			3573 => std_logic_vector(to_unsigned(75, 8)),
			3574 => std_logic_vector(to_unsigned(38, 8)),
			3575 => std_logic_vector(to_unsigned(199, 8)),
			3576 => std_logic_vector(to_unsigned(73, 8)),
			3577 => std_logic_vector(to_unsigned(210, 8)),
			3578 => std_logic_vector(to_unsigned(4, 8)),
			3579 => std_logic_vector(to_unsigned(29, 8)),
			3580 => std_logic_vector(to_unsigned(68, 8)),
			3581 => std_logic_vector(to_unsigned(74, 8)),
			3582 => std_logic_vector(to_unsigned(170, 8)),
			3583 => std_logic_vector(to_unsigned(13, 8)),
			3584 => std_logic_vector(to_unsigned(177, 8)),
			3585 => std_logic_vector(to_unsigned(36, 8)),
			3586 => std_logic_vector(to_unsigned(57, 8)),
			3587 => std_logic_vector(to_unsigned(147, 8)),
			3588 => std_logic_vector(to_unsigned(225, 8)),
			3589 => std_logic_vector(to_unsigned(13, 8)),
			3590 => std_logic_vector(to_unsigned(215, 8)),
			3591 => std_logic_vector(to_unsigned(254, 8)),
			3592 => std_logic_vector(to_unsigned(143, 8)),
			3593 => std_logic_vector(to_unsigned(241, 8)),
			3594 => std_logic_vector(to_unsigned(118, 8)),
			3595 => std_logic_vector(to_unsigned(2, 8)),
			3596 => std_logic_vector(to_unsigned(194, 8)),
			3597 => std_logic_vector(to_unsigned(141, 8)),
			3598 => std_logic_vector(to_unsigned(26, 8)),
			3599 => std_logic_vector(to_unsigned(159, 8)),
			3600 => std_logic_vector(to_unsigned(222, 8)),
			3601 => std_logic_vector(to_unsigned(131, 8)),
			3602 => std_logic_vector(to_unsigned(36, 8)),
			3603 => std_logic_vector(to_unsigned(53, 8)),
			3604 => std_logic_vector(to_unsigned(124, 8)),
			3605 => std_logic_vector(to_unsigned(85, 8)),
			3606 => std_logic_vector(to_unsigned(184, 8)),
			3607 => std_logic_vector(to_unsigned(36, 8)),
			3608 => std_logic_vector(to_unsigned(247, 8)),
			3609 => std_logic_vector(to_unsigned(236, 8)),
			3610 => std_logic_vector(to_unsigned(54, 8)),
			3611 => std_logic_vector(to_unsigned(119, 8)),
			others => (others => '0'));      

signal RAM2: ram_type := (0 => std_logic_vector(to_unsigned(69, 8)),
			1 => std_logic_vector(to_unsigned(24, 8)),
			2 => std_logic_vector(to_unsigned(128, 8)),
			3 => std_logic_vector(to_unsigned(52, 8)),
			4 => std_logic_vector(to_unsigned(241, 8)),
			5 => std_logic_vector(to_unsigned(188, 8)),
			6 => std_logic_vector(to_unsigned(70, 8)),
			7 => std_logic_vector(to_unsigned(128, 8)),
			8 => std_logic_vector(to_unsigned(71, 8)),
			9 => std_logic_vector(to_unsigned(118, 8)),
			10 => std_logic_vector(to_unsigned(30, 8)),
			11 => std_logic_vector(to_unsigned(172, 8)),
			12 => std_logic_vector(to_unsigned(227, 8)),
			13 => std_logic_vector(to_unsigned(79, 8)),
			14 => std_logic_vector(to_unsigned(40, 8)),
			15 => std_logic_vector(to_unsigned(117, 8)),
			16 => std_logic_vector(to_unsigned(49, 8)),
			17 => std_logic_vector(to_unsigned(79, 8)),
			18 => std_logic_vector(to_unsigned(193, 8)),
			19 => std_logic_vector(to_unsigned(19, 8)),
			20 => std_logic_vector(to_unsigned(28, 8)),
			21 => std_logic_vector(to_unsigned(199, 8)),
			22 => std_logic_vector(to_unsigned(119, 8)),
			23 => std_logic_vector(to_unsigned(210, 8)),
			24 => std_logic_vector(to_unsigned(143, 8)),
			25 => std_logic_vector(to_unsigned(238, 8)),
			26 => std_logic_vector(to_unsigned(27, 8)),
			27 => std_logic_vector(to_unsigned(255, 8)),
			28 => std_logic_vector(to_unsigned(155, 8)),
			29 => std_logic_vector(to_unsigned(147, 8)),
			30 => std_logic_vector(to_unsigned(169, 8)),
			31 => std_logic_vector(to_unsigned(153, 8)),
			32 => std_logic_vector(to_unsigned(204, 8)),
			33 => std_logic_vector(to_unsigned(234, 8)),
			34 => std_logic_vector(to_unsigned(3, 8)),
			35 => std_logic_vector(to_unsigned(5, 8)),
			36 => std_logic_vector(to_unsigned(65, 8)),
			37 => std_logic_vector(to_unsigned(44, 8)),
			38 => std_logic_vector(to_unsigned(228, 8)),
			39 => std_logic_vector(to_unsigned(93, 8)),
			40 => std_logic_vector(to_unsigned(8, 8)),
			41 => std_logic_vector(to_unsigned(93, 8)),
			42 => std_logic_vector(to_unsigned(30, 8)),
			43 => std_logic_vector(to_unsigned(119, 8)),
			44 => std_logic_vector(to_unsigned(114, 8)),
			45 => std_logic_vector(to_unsigned(84, 8)),
			46 => std_logic_vector(to_unsigned(13, 8)),
			47 => std_logic_vector(to_unsigned(84, 8)),
			48 => std_logic_vector(to_unsigned(247, 8)),
			49 => std_logic_vector(to_unsigned(99, 8)),
			50 => std_logic_vector(to_unsigned(217, 8)),
			51 => std_logic_vector(to_unsigned(204, 8)),
			52 => std_logic_vector(to_unsigned(252, 8)),
			53 => std_logic_vector(to_unsigned(2, 8)),
			54 => std_logic_vector(to_unsigned(99, 8)),
			55 => std_logic_vector(to_unsigned(176, 8)),
			56 => std_logic_vector(to_unsigned(40, 8)),
			57 => std_logic_vector(to_unsigned(255, 8)),
			58 => std_logic_vector(to_unsigned(96, 8)),
			59 => std_logic_vector(to_unsigned(171, 8)),
			60 => std_logic_vector(to_unsigned(90, 8)),
			61 => std_logic_vector(to_unsigned(231, 8)),
			62 => std_logic_vector(to_unsigned(32, 8)),
			63 => std_logic_vector(to_unsigned(25, 8)),
			64 => std_logic_vector(to_unsigned(12, 8)),
			65 => std_logic_vector(to_unsigned(150, 8)),
			66 => std_logic_vector(to_unsigned(21, 8)),
			67 => std_logic_vector(to_unsigned(85, 8)),
			68 => std_logic_vector(to_unsigned(21, 8)),
			69 => std_logic_vector(to_unsigned(39, 8)),
			70 => std_logic_vector(to_unsigned(59, 8)),
			71 => std_logic_vector(to_unsigned(61, 8)),
			72 => std_logic_vector(to_unsigned(45, 8)),
			73 => std_logic_vector(to_unsigned(109, 8)),
			74 => std_logic_vector(to_unsigned(11, 8)),
			75 => std_logic_vector(to_unsigned(16, 8)),
			76 => std_logic_vector(to_unsigned(183, 8)),
			77 => std_logic_vector(to_unsigned(177, 8)),
			78 => std_logic_vector(to_unsigned(227, 8)),
			79 => std_logic_vector(to_unsigned(15, 8)),
			80 => std_logic_vector(to_unsigned(123, 8)),
			81 => std_logic_vector(to_unsigned(95, 8)),
			82 => std_logic_vector(to_unsigned(134, 8)),
			83 => std_logic_vector(to_unsigned(56, 8)),
			84 => std_logic_vector(to_unsigned(6, 8)),
			85 => std_logic_vector(to_unsigned(206, 8)),
			86 => std_logic_vector(to_unsigned(94, 8)),
			87 => std_logic_vector(to_unsigned(8, 8)),
			88 => std_logic_vector(to_unsigned(81, 8)),
			89 => std_logic_vector(to_unsigned(15, 8)),
			90 => std_logic_vector(to_unsigned(61, 8)),
			91 => std_logic_vector(to_unsigned(24, 8)),
			92 => std_logic_vector(to_unsigned(173, 8)),
			93 => std_logic_vector(to_unsigned(188, 8)),
			94 => std_logic_vector(to_unsigned(229, 8)),
			95 => std_logic_vector(to_unsigned(161, 8)),
			96 => std_logic_vector(to_unsigned(204, 8)),
			97 => std_logic_vector(to_unsigned(34, 8)),
			98 => std_logic_vector(to_unsigned(6, 8)),
			99 => std_logic_vector(to_unsigned(167, 8)),
			100 => std_logic_vector(to_unsigned(174, 8)),
			101 => std_logic_vector(to_unsigned(23, 8)),
			102 => std_logic_vector(to_unsigned(203, 8)),
			103 => std_logic_vector(to_unsigned(108, 8)),
			104 => std_logic_vector(to_unsigned(148, 8)),
			105 => std_logic_vector(to_unsigned(176, 8)),
			106 => std_logic_vector(to_unsigned(148, 8)),
			107 => std_logic_vector(to_unsigned(183, 8)),
			108 => std_logic_vector(to_unsigned(37, 8)),
			109 => std_logic_vector(to_unsigned(52, 8)),
			110 => std_logic_vector(to_unsigned(196, 8)),
			111 => std_logic_vector(to_unsigned(44, 8)),
			112 => std_logic_vector(to_unsigned(238, 8)),
			113 => std_logic_vector(to_unsigned(142, 8)),
			114 => std_logic_vector(to_unsigned(239, 8)),
			115 => std_logic_vector(to_unsigned(119, 8)),
			116 => std_logic_vector(to_unsigned(185, 8)),
			117 => std_logic_vector(to_unsigned(35, 8)),
			118 => std_logic_vector(to_unsigned(42, 8)),
			119 => std_logic_vector(to_unsigned(171, 8)),
			120 => std_logic_vector(to_unsigned(252, 8)),
			121 => std_logic_vector(to_unsigned(31, 8)),
			122 => std_logic_vector(to_unsigned(137, 8)),
			123 => std_logic_vector(to_unsigned(60, 8)),
			124 => std_logic_vector(to_unsigned(92, 8)),
			125 => std_logic_vector(to_unsigned(9, 8)),
			126 => std_logic_vector(to_unsigned(247, 8)),
			127 => std_logic_vector(to_unsigned(26, 8)),
			128 => std_logic_vector(to_unsigned(244, 8)),
			129 => std_logic_vector(to_unsigned(58, 8)),
			130 => std_logic_vector(to_unsigned(217, 8)),
			131 => std_logic_vector(to_unsigned(44, 8)),
			132 => std_logic_vector(to_unsigned(142, 8)),
			133 => std_logic_vector(to_unsigned(196, 8)),
			134 => std_logic_vector(to_unsigned(89, 8)),
			135 => std_logic_vector(to_unsigned(63, 8)),
			136 => std_logic_vector(to_unsigned(41, 8)),
			137 => std_logic_vector(to_unsigned(253, 8)),
			138 => std_logic_vector(to_unsigned(251, 8)),
			139 => std_logic_vector(to_unsigned(253, 8)),
			140 => std_logic_vector(to_unsigned(181, 8)),
			141 => std_logic_vector(to_unsigned(184, 8)),
			142 => std_logic_vector(to_unsigned(194, 8)),
			143 => std_logic_vector(to_unsigned(66, 8)),
			144 => std_logic_vector(to_unsigned(187, 8)),
			145 => std_logic_vector(to_unsigned(11, 8)),
			146 => std_logic_vector(to_unsigned(70, 8)),
			147 => std_logic_vector(to_unsigned(168, 8)),
			148 => std_logic_vector(to_unsigned(44, 8)),
			149 => std_logic_vector(to_unsigned(146, 8)),
			150 => std_logic_vector(to_unsigned(172, 8)),
			151 => std_logic_vector(to_unsigned(221, 8)),
			152 => std_logic_vector(to_unsigned(244, 8)),
			153 => std_logic_vector(to_unsigned(93, 8)),
			154 => std_logic_vector(to_unsigned(1, 8)),
			155 => std_logic_vector(to_unsigned(82, 8)),
			156 => std_logic_vector(to_unsigned(129, 8)),
			157 => std_logic_vector(to_unsigned(173, 8)),
			158 => std_logic_vector(to_unsigned(69, 8)),
			159 => std_logic_vector(to_unsigned(51, 8)),
			160 => std_logic_vector(to_unsigned(92, 8)),
			161 => std_logic_vector(to_unsigned(175, 8)),
			162 => std_logic_vector(to_unsigned(186, 8)),
			163 => std_logic_vector(to_unsigned(164, 8)),
			164 => std_logic_vector(to_unsigned(233, 8)),
			165 => std_logic_vector(to_unsigned(120, 8)),
			166 => std_logic_vector(to_unsigned(30, 8)),
			167 => std_logic_vector(to_unsigned(105, 8)),
			168 => std_logic_vector(to_unsigned(246, 8)),
			169 => std_logic_vector(to_unsigned(215, 8)),
			170 => std_logic_vector(to_unsigned(238, 8)),
			171 => std_logic_vector(to_unsigned(57, 8)),
			172 => std_logic_vector(to_unsigned(146, 8)),
			173 => std_logic_vector(to_unsigned(245, 8)),
			174 => std_logic_vector(to_unsigned(142, 8)),
			175 => std_logic_vector(to_unsigned(94, 8)),
			176 => std_logic_vector(to_unsigned(197, 8)),
			177 => std_logic_vector(to_unsigned(75, 8)),
			178 => std_logic_vector(to_unsigned(23, 8)),
			179 => std_logic_vector(to_unsigned(204, 8)),
			180 => std_logic_vector(to_unsigned(99, 8)),
			181 => std_logic_vector(to_unsigned(172, 8)),
			182 => std_logic_vector(to_unsigned(135, 8)),
			183 => std_logic_vector(to_unsigned(31, 8)),
			184 => std_logic_vector(to_unsigned(73, 8)),
			185 => std_logic_vector(to_unsigned(189, 8)),
			186 => std_logic_vector(to_unsigned(35, 8)),
			187 => std_logic_vector(to_unsigned(97, 8)),
			188 => std_logic_vector(to_unsigned(175, 8)),
			189 => std_logic_vector(to_unsigned(219, 8)),
			190 => std_logic_vector(to_unsigned(37, 8)),
			191 => std_logic_vector(to_unsigned(102, 8)),
			192 => std_logic_vector(to_unsigned(107, 8)),
			193 => std_logic_vector(to_unsigned(124, 8)),
			194 => std_logic_vector(to_unsigned(34, 8)),
			195 => std_logic_vector(to_unsigned(82, 8)),
			196 => std_logic_vector(to_unsigned(206, 8)),
			197 => std_logic_vector(to_unsigned(105, 8)),
			198 => std_logic_vector(to_unsigned(151, 8)),
			199 => std_logic_vector(to_unsigned(46, 8)),
			200 => std_logic_vector(to_unsigned(94, 8)),
			201 => std_logic_vector(to_unsigned(180, 8)),
			202 => std_logic_vector(to_unsigned(42, 8)),
			203 => std_logic_vector(to_unsigned(136, 8)),
			204 => std_logic_vector(to_unsigned(245, 8)),
			205 => std_logic_vector(to_unsigned(103, 8)),
			206 => std_logic_vector(to_unsigned(127, 8)),
			207 => std_logic_vector(to_unsigned(181, 8)),
			208 => std_logic_vector(to_unsigned(128, 8)),
			209 => std_logic_vector(to_unsigned(234, 8)),
			210 => std_logic_vector(to_unsigned(89, 8)),
			211 => std_logic_vector(to_unsigned(255, 8)),
			212 => std_logic_vector(to_unsigned(123, 8)),
			213 => std_logic_vector(to_unsigned(183, 8)),
			214 => std_logic_vector(to_unsigned(104, 8)),
			215 => std_logic_vector(to_unsigned(90, 8)),
			216 => std_logic_vector(to_unsigned(2, 8)),
			217 => std_logic_vector(to_unsigned(143, 8)),
			218 => std_logic_vector(to_unsigned(200, 8)),
			219 => std_logic_vector(to_unsigned(242, 8)),
			220 => std_logic_vector(to_unsigned(166, 8)),
			221 => std_logic_vector(to_unsigned(112, 8)),
			222 => std_logic_vector(to_unsigned(150, 8)),
			223 => std_logic_vector(to_unsigned(11, 8)),
			224 => std_logic_vector(to_unsigned(158, 8)),
			225 => std_logic_vector(to_unsigned(92, 8)),
			226 => std_logic_vector(to_unsigned(88, 8)),
			227 => std_logic_vector(to_unsigned(216, 8)),
			228 => std_logic_vector(to_unsigned(86, 8)),
			229 => std_logic_vector(to_unsigned(177, 8)),
			230 => std_logic_vector(to_unsigned(96, 8)),
			231 => std_logic_vector(to_unsigned(232, 8)),
			232 => std_logic_vector(to_unsigned(153, 8)),
			233 => std_logic_vector(to_unsigned(194, 8)),
			234 => std_logic_vector(to_unsigned(243, 8)),
			235 => std_logic_vector(to_unsigned(14, 8)),
			236 => std_logic_vector(to_unsigned(41, 8)),
			237 => std_logic_vector(to_unsigned(198, 8)),
			238 => std_logic_vector(to_unsigned(118, 8)),
			239 => std_logic_vector(to_unsigned(14, 8)),
			240 => std_logic_vector(to_unsigned(107, 8)),
			241 => std_logic_vector(to_unsigned(169, 8)),
			242 => std_logic_vector(to_unsigned(125, 8)),
			243 => std_logic_vector(to_unsigned(156, 8)),
			244 => std_logic_vector(to_unsigned(93, 8)),
			245 => std_logic_vector(to_unsigned(88, 8)),
			246 => std_logic_vector(to_unsigned(84, 8)),
			247 => std_logic_vector(to_unsigned(147, 8)),
			248 => std_logic_vector(to_unsigned(240, 8)),
			249 => std_logic_vector(to_unsigned(220, 8)),
			250 => std_logic_vector(to_unsigned(71, 8)),
			251 => std_logic_vector(to_unsigned(44, 8)),
			252 => std_logic_vector(to_unsigned(171, 8)),
			253 => std_logic_vector(to_unsigned(59, 8)),
			254 => std_logic_vector(to_unsigned(204, 8)),
			255 => std_logic_vector(to_unsigned(193, 8)),
			256 => std_logic_vector(to_unsigned(27, 8)),
			257 => std_logic_vector(to_unsigned(131, 8)),
			258 => std_logic_vector(to_unsigned(142, 8)),
			259 => std_logic_vector(to_unsigned(150, 8)),
			260 => std_logic_vector(to_unsigned(158, 8)),
			261 => std_logic_vector(to_unsigned(105, 8)),
			262 => std_logic_vector(to_unsigned(65, 8)),
			263 => std_logic_vector(to_unsigned(187, 8)),
			264 => std_logic_vector(to_unsigned(210, 8)),
			265 => std_logic_vector(to_unsigned(80, 8)),
			266 => std_logic_vector(to_unsigned(83, 8)),
			267 => std_logic_vector(to_unsigned(254, 8)),
			268 => std_logic_vector(to_unsigned(168, 8)),
			269 => std_logic_vector(to_unsigned(200, 8)),
			270 => std_logic_vector(to_unsigned(87, 8)),
			271 => std_logic_vector(to_unsigned(95, 8)),
			272 => std_logic_vector(to_unsigned(60, 8)),
			273 => std_logic_vector(to_unsigned(244, 8)),
			274 => std_logic_vector(to_unsigned(11, 8)),
			275 => std_logic_vector(to_unsigned(55, 8)),
			276 => std_logic_vector(to_unsigned(110, 8)),
			277 => std_logic_vector(to_unsigned(61, 8)),
			278 => std_logic_vector(to_unsigned(254, 8)),
			279 => std_logic_vector(to_unsigned(13, 8)),
			280 => std_logic_vector(to_unsigned(166, 8)),
			281 => std_logic_vector(to_unsigned(82, 8)),
			282 => std_logic_vector(to_unsigned(13, 8)),
			283 => std_logic_vector(to_unsigned(23, 8)),
			284 => std_logic_vector(to_unsigned(62, 8)),
			285 => std_logic_vector(to_unsigned(216, 8)),
			286 => std_logic_vector(to_unsigned(63, 8)),
			287 => std_logic_vector(to_unsigned(244, 8)),
			288 => std_logic_vector(to_unsigned(37, 8)),
			289 => std_logic_vector(to_unsigned(253, 8)),
			290 => std_logic_vector(to_unsigned(210, 8)),
			291 => std_logic_vector(to_unsigned(199, 8)),
			292 => std_logic_vector(to_unsigned(186, 8)),
			293 => std_logic_vector(to_unsigned(50, 8)),
			294 => std_logic_vector(to_unsigned(188, 8)),
			295 => std_logic_vector(to_unsigned(79, 8)),
			296 => std_logic_vector(to_unsigned(122, 8)),
			297 => std_logic_vector(to_unsigned(202, 8)),
			298 => std_logic_vector(to_unsigned(223, 8)),
			299 => std_logic_vector(to_unsigned(217, 8)),
			300 => std_logic_vector(to_unsigned(171, 8)),
			301 => std_logic_vector(to_unsigned(231, 8)),
			302 => std_logic_vector(to_unsigned(134, 8)),
			303 => std_logic_vector(to_unsigned(24, 8)),
			304 => std_logic_vector(to_unsigned(79, 8)),
			305 => std_logic_vector(to_unsigned(119, 8)),
			306 => std_logic_vector(to_unsigned(125, 8)),
			307 => std_logic_vector(to_unsigned(10, 8)),
			308 => std_logic_vector(to_unsigned(99, 8)),
			309 => std_logic_vector(to_unsigned(203, 8)),
			310 => std_logic_vector(to_unsigned(160, 8)),
			311 => std_logic_vector(to_unsigned(125, 8)),
			312 => std_logic_vector(to_unsigned(30, 8)),
			313 => std_logic_vector(to_unsigned(213, 8)),
			314 => std_logic_vector(to_unsigned(33, 8)),
			315 => std_logic_vector(to_unsigned(17, 8)),
			316 => std_logic_vector(to_unsigned(132, 8)),
			317 => std_logic_vector(to_unsigned(71, 8)),
			318 => std_logic_vector(to_unsigned(111, 8)),
			319 => std_logic_vector(to_unsigned(22, 8)),
			320 => std_logic_vector(to_unsigned(58, 8)),
			321 => std_logic_vector(to_unsigned(194, 8)),
			322 => std_logic_vector(to_unsigned(54, 8)),
			323 => std_logic_vector(to_unsigned(78, 8)),
			324 => std_logic_vector(to_unsigned(42, 8)),
			325 => std_logic_vector(to_unsigned(45, 8)),
			326 => std_logic_vector(to_unsigned(99, 8)),
			327 => std_logic_vector(to_unsigned(155, 8)),
			328 => std_logic_vector(to_unsigned(153, 8)),
			329 => std_logic_vector(to_unsigned(173, 8)),
			330 => std_logic_vector(to_unsigned(7, 8)),
			331 => std_logic_vector(to_unsigned(220, 8)),
			332 => std_logic_vector(to_unsigned(136, 8)),
			333 => std_logic_vector(to_unsigned(162, 8)),
			334 => std_logic_vector(to_unsigned(61, 8)),
			335 => std_logic_vector(to_unsigned(194, 8)),
			336 => std_logic_vector(to_unsigned(104, 8)),
			337 => std_logic_vector(to_unsigned(253, 8)),
			338 => std_logic_vector(to_unsigned(221, 8)),
			339 => std_logic_vector(to_unsigned(173, 8)),
			340 => std_logic_vector(to_unsigned(212, 8)),
			341 => std_logic_vector(to_unsigned(28, 8)),
			342 => std_logic_vector(to_unsigned(170, 8)),
			343 => std_logic_vector(to_unsigned(59, 8)),
			344 => std_logic_vector(to_unsigned(147, 8)),
			345 => std_logic_vector(to_unsigned(8, 8)),
			346 => std_logic_vector(to_unsigned(235, 8)),
			347 => std_logic_vector(to_unsigned(118, 8)),
			348 => std_logic_vector(to_unsigned(117, 8)),
			349 => std_logic_vector(to_unsigned(189, 8)),
			350 => std_logic_vector(to_unsigned(115, 8)),
			351 => std_logic_vector(to_unsigned(202, 8)),
			352 => std_logic_vector(to_unsigned(228, 8)),
			353 => std_logic_vector(to_unsigned(153, 8)),
			354 => std_logic_vector(to_unsigned(87, 8)),
			355 => std_logic_vector(to_unsigned(57, 8)),
			356 => std_logic_vector(to_unsigned(74, 8)),
			357 => std_logic_vector(to_unsigned(212, 8)),
			358 => std_logic_vector(to_unsigned(127, 8)),
			359 => std_logic_vector(to_unsigned(19, 8)),
			360 => std_logic_vector(to_unsigned(181, 8)),
			361 => std_logic_vector(to_unsigned(135, 8)),
			362 => std_logic_vector(to_unsigned(122, 8)),
			363 => std_logic_vector(to_unsigned(110, 8)),
			364 => std_logic_vector(to_unsigned(7, 8)),
			365 => std_logic_vector(to_unsigned(134, 8)),
			366 => std_logic_vector(to_unsigned(6, 8)),
			367 => std_logic_vector(to_unsigned(85, 8)),
			368 => std_logic_vector(to_unsigned(29, 8)),
			369 => std_logic_vector(to_unsigned(19, 8)),
			370 => std_logic_vector(to_unsigned(34, 8)),
			371 => std_logic_vector(to_unsigned(139, 8)),
			372 => std_logic_vector(to_unsigned(30, 8)),
			373 => std_logic_vector(to_unsigned(86, 8)),
			374 => std_logic_vector(to_unsigned(3, 8)),
			375 => std_logic_vector(to_unsigned(132, 8)),
			376 => std_logic_vector(to_unsigned(5, 8)),
			377 => std_logic_vector(to_unsigned(115, 8)),
			378 => std_logic_vector(to_unsigned(143, 8)),
			379 => std_logic_vector(to_unsigned(6, 8)),
			380 => std_logic_vector(to_unsigned(224, 8)),
			381 => std_logic_vector(to_unsigned(208, 8)),
			382 => std_logic_vector(to_unsigned(36, 8)),
			383 => std_logic_vector(to_unsigned(25, 8)),
			384 => std_logic_vector(to_unsigned(42, 8)),
			385 => std_logic_vector(to_unsigned(152, 8)),
			386 => std_logic_vector(to_unsigned(18, 8)),
			387 => std_logic_vector(to_unsigned(31, 8)),
			388 => std_logic_vector(to_unsigned(132, 8)),
			389 => std_logic_vector(to_unsigned(145, 8)),
			390 => std_logic_vector(to_unsigned(199, 8)),
			391 => std_logic_vector(to_unsigned(48, 8)),
			392 => std_logic_vector(to_unsigned(119, 8)),
			393 => std_logic_vector(to_unsigned(108, 8)),
			394 => std_logic_vector(to_unsigned(27, 8)),
			395 => std_logic_vector(to_unsigned(235, 8)),
			396 => std_logic_vector(to_unsigned(112, 8)),
			397 => std_logic_vector(to_unsigned(112, 8)),
			398 => std_logic_vector(to_unsigned(238, 8)),
			399 => std_logic_vector(to_unsigned(184, 8)),
			400 => std_logic_vector(to_unsigned(179, 8)),
			401 => std_logic_vector(to_unsigned(106, 8)),
			402 => std_logic_vector(to_unsigned(95, 8)),
			403 => std_logic_vector(to_unsigned(10, 8)),
			404 => std_logic_vector(to_unsigned(226, 8)),
			405 => std_logic_vector(to_unsigned(250, 8)),
			406 => std_logic_vector(to_unsigned(223, 8)),
			407 => std_logic_vector(to_unsigned(44, 8)),
			408 => std_logic_vector(to_unsigned(98, 8)),
			409 => std_logic_vector(to_unsigned(255, 8)),
			410 => std_logic_vector(to_unsigned(191, 8)),
			411 => std_logic_vector(to_unsigned(216, 8)),
			412 => std_logic_vector(to_unsigned(234, 8)),
			413 => std_logic_vector(to_unsigned(52, 8)),
			414 => std_logic_vector(to_unsigned(154, 8)),
			415 => std_logic_vector(to_unsigned(57, 8)),
			416 => std_logic_vector(to_unsigned(58, 8)),
			417 => std_logic_vector(to_unsigned(106, 8)),
			418 => std_logic_vector(to_unsigned(132, 8)),
			419 => std_logic_vector(to_unsigned(101, 8)),
			420 => std_logic_vector(to_unsigned(213, 8)),
			421 => std_logic_vector(to_unsigned(202, 8)),
			422 => std_logic_vector(to_unsigned(209, 8)),
			423 => std_logic_vector(to_unsigned(188, 8)),
			424 => std_logic_vector(to_unsigned(142, 8)),
			425 => std_logic_vector(to_unsigned(25, 8)),
			426 => std_logic_vector(to_unsigned(111, 8)),
			427 => std_logic_vector(to_unsigned(200, 8)),
			428 => std_logic_vector(to_unsigned(40, 8)),
			429 => std_logic_vector(to_unsigned(247, 8)),
			430 => std_logic_vector(to_unsigned(52, 8)),
			431 => std_logic_vector(to_unsigned(176, 8)),
			432 => std_logic_vector(to_unsigned(83, 8)),
			433 => std_logic_vector(to_unsigned(173, 8)),
			434 => std_logic_vector(to_unsigned(224, 8)),
			435 => std_logic_vector(to_unsigned(96, 8)),
			436 => std_logic_vector(to_unsigned(193, 8)),
			437 => std_logic_vector(to_unsigned(134, 8)),
			438 => std_logic_vector(to_unsigned(95, 8)),
			439 => std_logic_vector(to_unsigned(52, 8)),
			440 => std_logic_vector(to_unsigned(102, 8)),
			441 => std_logic_vector(to_unsigned(1, 8)),
			442 => std_logic_vector(to_unsigned(113, 8)),
			443 => std_logic_vector(to_unsigned(41, 8)),
			444 => std_logic_vector(to_unsigned(58, 8)),
			445 => std_logic_vector(to_unsigned(15, 8)),
			446 => std_logic_vector(to_unsigned(85, 8)),
			447 => std_logic_vector(to_unsigned(154, 8)),
			448 => std_logic_vector(to_unsigned(98, 8)),
			449 => std_logic_vector(to_unsigned(56, 8)),
			450 => std_logic_vector(to_unsigned(23, 8)),
			451 => std_logic_vector(to_unsigned(227, 8)),
			452 => std_logic_vector(to_unsigned(34, 8)),
			453 => std_logic_vector(to_unsigned(9, 8)),
			454 => std_logic_vector(to_unsigned(127, 8)),
			455 => std_logic_vector(to_unsigned(154, 8)),
			456 => std_logic_vector(to_unsigned(171, 8)),
			457 => std_logic_vector(to_unsigned(75, 8)),
			458 => std_logic_vector(to_unsigned(48, 8)),
			459 => std_logic_vector(to_unsigned(211, 8)),
			460 => std_logic_vector(to_unsigned(205, 8)),
			461 => std_logic_vector(to_unsigned(6, 8)),
			462 => std_logic_vector(to_unsigned(195, 8)),
			463 => std_logic_vector(to_unsigned(34, 8)),
			464 => std_logic_vector(to_unsigned(119, 8)),
			465 => std_logic_vector(to_unsigned(68, 8)),
			466 => std_logic_vector(to_unsigned(17, 8)),
			467 => std_logic_vector(to_unsigned(160, 8)),
			468 => std_logic_vector(to_unsigned(11, 8)),
			469 => std_logic_vector(to_unsigned(17, 8)),
			470 => std_logic_vector(to_unsigned(91, 8)),
			471 => std_logic_vector(to_unsigned(108, 8)),
			472 => std_logic_vector(to_unsigned(7, 8)),
			473 => std_logic_vector(to_unsigned(43, 8)),
			474 => std_logic_vector(to_unsigned(234, 8)),
			475 => std_logic_vector(to_unsigned(18, 8)),
			476 => std_logic_vector(to_unsigned(96, 8)),
			477 => std_logic_vector(to_unsigned(47, 8)),
			478 => std_logic_vector(to_unsigned(243, 8)),
			479 => std_logic_vector(to_unsigned(245, 8)),
			480 => std_logic_vector(to_unsigned(201, 8)),
			481 => std_logic_vector(to_unsigned(128, 8)),
			482 => std_logic_vector(to_unsigned(39, 8)),
			483 => std_logic_vector(to_unsigned(59, 8)),
			484 => std_logic_vector(to_unsigned(54, 8)),
			485 => std_logic_vector(to_unsigned(135, 8)),
			486 => std_logic_vector(to_unsigned(7, 8)),
			487 => std_logic_vector(to_unsigned(60, 8)),
			488 => std_logic_vector(to_unsigned(91, 8)),
			489 => std_logic_vector(to_unsigned(243, 8)),
			490 => std_logic_vector(to_unsigned(236, 8)),
			491 => std_logic_vector(to_unsigned(75, 8)),
			492 => std_logic_vector(to_unsigned(157, 8)),
			493 => std_logic_vector(to_unsigned(147, 8)),
			494 => std_logic_vector(to_unsigned(142, 8)),
			495 => std_logic_vector(to_unsigned(16, 8)),
			496 => std_logic_vector(to_unsigned(238, 8)),
			497 => std_logic_vector(to_unsigned(53, 8)),
			498 => std_logic_vector(to_unsigned(108, 8)),
			499 => std_logic_vector(to_unsigned(204, 8)),
			500 => std_logic_vector(to_unsigned(64, 8)),
			501 => std_logic_vector(to_unsigned(195, 8)),
			502 => std_logic_vector(to_unsigned(114, 8)),
			503 => std_logic_vector(to_unsigned(124, 8)),
			504 => std_logic_vector(to_unsigned(198, 8)),
			505 => std_logic_vector(to_unsigned(10, 8)),
			506 => std_logic_vector(to_unsigned(249, 8)),
			507 => std_logic_vector(to_unsigned(168, 8)),
			508 => std_logic_vector(to_unsigned(83, 8)),
			509 => std_logic_vector(to_unsigned(169, 8)),
			510 => std_logic_vector(to_unsigned(228, 8)),
			511 => std_logic_vector(to_unsigned(127, 8)),
			512 => std_logic_vector(to_unsigned(217, 8)),
			513 => std_logic_vector(to_unsigned(239, 8)),
			514 => std_logic_vector(to_unsigned(80, 8)),
			515 => std_logic_vector(to_unsigned(185, 8)),
			516 => std_logic_vector(to_unsigned(160, 8)),
			517 => std_logic_vector(to_unsigned(234, 8)),
			518 => std_logic_vector(to_unsigned(159, 8)),
			519 => std_logic_vector(to_unsigned(92, 8)),
			520 => std_logic_vector(to_unsigned(106, 8)),
			521 => std_logic_vector(to_unsigned(190, 8)),
			522 => std_logic_vector(to_unsigned(232, 8)),
			523 => std_logic_vector(to_unsigned(122, 8)),
			524 => std_logic_vector(to_unsigned(131, 8)),
			525 => std_logic_vector(to_unsigned(178, 8)),
			526 => std_logic_vector(to_unsigned(164, 8)),
			527 => std_logic_vector(to_unsigned(161, 8)),
			528 => std_logic_vector(to_unsigned(210, 8)),
			529 => std_logic_vector(to_unsigned(226, 8)),
			530 => std_logic_vector(to_unsigned(160, 8)),
			531 => std_logic_vector(to_unsigned(72, 8)),
			532 => std_logic_vector(to_unsigned(22, 8)),
			533 => std_logic_vector(to_unsigned(1, 8)),
			534 => std_logic_vector(to_unsigned(44, 8)),
			535 => std_logic_vector(to_unsigned(146, 8)),
			536 => std_logic_vector(to_unsigned(217, 8)),
			537 => std_logic_vector(to_unsigned(177, 8)),
			538 => std_logic_vector(to_unsigned(109, 8)),
			539 => std_logic_vector(to_unsigned(191, 8)),
			540 => std_logic_vector(to_unsigned(133, 8)),
			541 => std_logic_vector(to_unsigned(157, 8)),
			542 => std_logic_vector(to_unsigned(106, 8)),
			543 => std_logic_vector(to_unsigned(118, 8)),
			544 => std_logic_vector(to_unsigned(9, 8)),
			545 => std_logic_vector(to_unsigned(7, 8)),
			546 => std_logic_vector(to_unsigned(94, 8)),
			547 => std_logic_vector(to_unsigned(172, 8)),
			548 => std_logic_vector(to_unsigned(115, 8)),
			549 => std_logic_vector(to_unsigned(220, 8)),
			550 => std_logic_vector(to_unsigned(192, 8)),
			551 => std_logic_vector(to_unsigned(197, 8)),
			552 => std_logic_vector(to_unsigned(216, 8)),
			553 => std_logic_vector(to_unsigned(24, 8)),
			554 => std_logic_vector(to_unsigned(225, 8)),
			555 => std_logic_vector(to_unsigned(61, 8)),
			556 => std_logic_vector(to_unsigned(104, 8)),
			557 => std_logic_vector(to_unsigned(121, 8)),
			558 => std_logic_vector(to_unsigned(207, 8)),
			559 => std_logic_vector(to_unsigned(251, 8)),
			560 => std_logic_vector(to_unsigned(141, 8)),
			561 => std_logic_vector(to_unsigned(111, 8)),
			562 => std_logic_vector(to_unsigned(27, 8)),
			563 => std_logic_vector(to_unsigned(142, 8)),
			564 => std_logic_vector(to_unsigned(238, 8)),
			565 => std_logic_vector(to_unsigned(56, 8)),
			566 => std_logic_vector(to_unsigned(45, 8)),
			567 => std_logic_vector(to_unsigned(70, 8)),
			568 => std_logic_vector(to_unsigned(6, 8)),
			569 => std_logic_vector(to_unsigned(162, 8)),
			570 => std_logic_vector(to_unsigned(207, 8)),
			571 => std_logic_vector(to_unsigned(142, 8)),
			572 => std_logic_vector(to_unsigned(79, 8)),
			573 => std_logic_vector(to_unsigned(188, 8)),
			574 => std_logic_vector(to_unsigned(183, 8)),
			575 => std_logic_vector(to_unsigned(162, 8)),
			576 => std_logic_vector(to_unsigned(168, 8)),
			577 => std_logic_vector(to_unsigned(183, 8)),
			578 => std_logic_vector(to_unsigned(11, 8)),
			579 => std_logic_vector(to_unsigned(235, 8)),
			580 => std_logic_vector(to_unsigned(0, 8)),
			581 => std_logic_vector(to_unsigned(58, 8)),
			582 => std_logic_vector(to_unsigned(235, 8)),
			583 => std_logic_vector(to_unsigned(219, 8)),
			584 => std_logic_vector(to_unsigned(248, 8)),
			585 => std_logic_vector(to_unsigned(177, 8)),
			586 => std_logic_vector(to_unsigned(115, 8)),
			587 => std_logic_vector(to_unsigned(187, 8)),
			588 => std_logic_vector(to_unsigned(224, 8)),
			589 => std_logic_vector(to_unsigned(86, 8)),
			590 => std_logic_vector(to_unsigned(160, 8)),
			591 => std_logic_vector(to_unsigned(41, 8)),
			592 => std_logic_vector(to_unsigned(219, 8)),
			593 => std_logic_vector(to_unsigned(198, 8)),
			594 => std_logic_vector(to_unsigned(183, 8)),
			595 => std_logic_vector(to_unsigned(49, 8)),
			596 => std_logic_vector(to_unsigned(223, 8)),
			597 => std_logic_vector(to_unsigned(151, 8)),
			598 => std_logic_vector(to_unsigned(151, 8)),
			599 => std_logic_vector(to_unsigned(215, 8)),
			600 => std_logic_vector(to_unsigned(139, 8)),
			601 => std_logic_vector(to_unsigned(134, 8)),
			602 => std_logic_vector(to_unsigned(233, 8)),
			603 => std_logic_vector(to_unsigned(176, 8)),
			604 => std_logic_vector(to_unsigned(35, 8)),
			605 => std_logic_vector(to_unsigned(153, 8)),
			606 => std_logic_vector(to_unsigned(97, 8)),
			607 => std_logic_vector(to_unsigned(208, 8)),
			608 => std_logic_vector(to_unsigned(216, 8)),
			609 => std_logic_vector(to_unsigned(92, 8)),
			610 => std_logic_vector(to_unsigned(120, 8)),
			611 => std_logic_vector(to_unsigned(25, 8)),
			612 => std_logic_vector(to_unsigned(215, 8)),
			613 => std_logic_vector(to_unsigned(235, 8)),
			614 => std_logic_vector(to_unsigned(208, 8)),
			615 => std_logic_vector(to_unsigned(245, 8)),
			616 => std_logic_vector(to_unsigned(17, 8)),
			617 => std_logic_vector(to_unsigned(222, 8)),
			618 => std_logic_vector(to_unsigned(173, 8)),
			619 => std_logic_vector(to_unsigned(0, 8)),
			620 => std_logic_vector(to_unsigned(188, 8)),
			621 => std_logic_vector(to_unsigned(201, 8)),
			622 => std_logic_vector(to_unsigned(103, 8)),
			623 => std_logic_vector(to_unsigned(103, 8)),
			624 => std_logic_vector(to_unsigned(79, 8)),
			625 => std_logic_vector(to_unsigned(232, 8)),
			626 => std_logic_vector(to_unsigned(170, 8)),
			627 => std_logic_vector(to_unsigned(241, 8)),
			628 => std_logic_vector(to_unsigned(243, 8)),
			629 => std_logic_vector(to_unsigned(160, 8)),
			630 => std_logic_vector(to_unsigned(158, 8)),
			631 => std_logic_vector(to_unsigned(166, 8)),
			632 => std_logic_vector(to_unsigned(84, 8)),
			633 => std_logic_vector(to_unsigned(137, 8)),
			634 => std_logic_vector(to_unsigned(57, 8)),
			635 => std_logic_vector(to_unsigned(29, 8)),
			636 => std_logic_vector(to_unsigned(10, 8)),
			637 => std_logic_vector(to_unsigned(36, 8)),
			638 => std_logic_vector(to_unsigned(226, 8)),
			639 => std_logic_vector(to_unsigned(91, 8)),
			640 => std_logic_vector(to_unsigned(170, 8)),
			641 => std_logic_vector(to_unsigned(212, 8)),
			642 => std_logic_vector(to_unsigned(169, 8)),
			643 => std_logic_vector(to_unsigned(132, 8)),
			644 => std_logic_vector(to_unsigned(112, 8)),
			645 => std_logic_vector(to_unsigned(246, 8)),
			646 => std_logic_vector(to_unsigned(235, 8)),
			647 => std_logic_vector(to_unsigned(197, 8)),
			648 => std_logic_vector(to_unsigned(249, 8)),
			649 => std_logic_vector(to_unsigned(61, 8)),
			650 => std_logic_vector(to_unsigned(57, 8)),
			651 => std_logic_vector(to_unsigned(146, 8)),
			652 => std_logic_vector(to_unsigned(79, 8)),
			653 => std_logic_vector(to_unsigned(122, 8)),
			654 => std_logic_vector(to_unsigned(116, 8)),
			655 => std_logic_vector(to_unsigned(159, 8)),
			656 => std_logic_vector(to_unsigned(173, 8)),
			657 => std_logic_vector(to_unsigned(1, 8)),
			658 => std_logic_vector(to_unsigned(4, 8)),
			659 => std_logic_vector(to_unsigned(71, 8)),
			660 => std_logic_vector(to_unsigned(205, 8)),
			661 => std_logic_vector(to_unsigned(81, 8)),
			662 => std_logic_vector(to_unsigned(95, 8)),
			663 => std_logic_vector(to_unsigned(35, 8)),
			664 => std_logic_vector(to_unsigned(241, 8)),
			665 => std_logic_vector(to_unsigned(20, 8)),
			666 => std_logic_vector(to_unsigned(49, 8)),
			667 => std_logic_vector(to_unsigned(3, 8)),
			668 => std_logic_vector(to_unsigned(121, 8)),
			669 => std_logic_vector(to_unsigned(188, 8)),
			670 => std_logic_vector(to_unsigned(197, 8)),
			671 => std_logic_vector(to_unsigned(17, 8)),
			672 => std_logic_vector(to_unsigned(44, 8)),
			673 => std_logic_vector(to_unsigned(228, 8)),
			674 => std_logic_vector(to_unsigned(142, 8)),
			675 => std_logic_vector(to_unsigned(10, 8)),
			676 => std_logic_vector(to_unsigned(235, 8)),
			677 => std_logic_vector(to_unsigned(8, 8)),
			678 => std_logic_vector(to_unsigned(88, 8)),
			679 => std_logic_vector(to_unsigned(98, 8)),
			680 => std_logic_vector(to_unsigned(24, 8)),
			681 => std_logic_vector(to_unsigned(47, 8)),
			682 => std_logic_vector(to_unsigned(201, 8)),
			683 => std_logic_vector(to_unsigned(221, 8)),
			684 => std_logic_vector(to_unsigned(136, 8)),
			685 => std_logic_vector(to_unsigned(145, 8)),
			686 => std_logic_vector(to_unsigned(76, 8)),
			687 => std_logic_vector(to_unsigned(241, 8)),
			688 => std_logic_vector(to_unsigned(206, 8)),
			689 => std_logic_vector(to_unsigned(214, 8)),
			690 => std_logic_vector(to_unsigned(43, 8)),
			691 => std_logic_vector(to_unsigned(93, 8)),
			692 => std_logic_vector(to_unsigned(235, 8)),
			693 => std_logic_vector(to_unsigned(85, 8)),
			694 => std_logic_vector(to_unsigned(217, 8)),
			695 => std_logic_vector(to_unsigned(139, 8)),
			696 => std_logic_vector(to_unsigned(207, 8)),
			697 => std_logic_vector(to_unsigned(173, 8)),
			698 => std_logic_vector(to_unsigned(115, 8)),
			699 => std_logic_vector(to_unsigned(113, 8)),
			700 => std_logic_vector(to_unsigned(222, 8)),
			701 => std_logic_vector(to_unsigned(219, 8)),
			702 => std_logic_vector(to_unsigned(99, 8)),
			703 => std_logic_vector(to_unsigned(55, 8)),
			704 => std_logic_vector(to_unsigned(181, 8)),
			705 => std_logic_vector(to_unsigned(182, 8)),
			706 => std_logic_vector(to_unsigned(127, 8)),
			707 => std_logic_vector(to_unsigned(19, 8)),
			708 => std_logic_vector(to_unsigned(73, 8)),
			709 => std_logic_vector(to_unsigned(56, 8)),
			710 => std_logic_vector(to_unsigned(50, 8)),
			711 => std_logic_vector(to_unsigned(234, 8)),
			712 => std_logic_vector(to_unsigned(67, 8)),
			713 => std_logic_vector(to_unsigned(125, 8)),
			714 => std_logic_vector(to_unsigned(11, 8)),
			715 => std_logic_vector(to_unsigned(131, 8)),
			716 => std_logic_vector(to_unsigned(148, 8)),
			717 => std_logic_vector(to_unsigned(94, 8)),
			718 => std_logic_vector(to_unsigned(218, 8)),
			719 => std_logic_vector(to_unsigned(42, 8)),
			720 => std_logic_vector(to_unsigned(245, 8)),
			721 => std_logic_vector(to_unsigned(192, 8)),
			722 => std_logic_vector(to_unsigned(101, 8)),
			723 => std_logic_vector(to_unsigned(243, 8)),
			724 => std_logic_vector(to_unsigned(92, 8)),
			725 => std_logic_vector(to_unsigned(171, 8)),
			726 => std_logic_vector(to_unsigned(91, 8)),
			727 => std_logic_vector(to_unsigned(148, 8)),
			728 => std_logic_vector(to_unsigned(43, 8)),
			729 => std_logic_vector(to_unsigned(125, 8)),
			730 => std_logic_vector(to_unsigned(146, 8)),
			731 => std_logic_vector(to_unsigned(229, 8)),
			732 => std_logic_vector(to_unsigned(160, 8)),
			733 => std_logic_vector(to_unsigned(236, 8)),
			734 => std_logic_vector(to_unsigned(173, 8)),
			735 => std_logic_vector(to_unsigned(84, 8)),
			736 => std_logic_vector(to_unsigned(223, 8)),
			737 => std_logic_vector(to_unsigned(51, 8)),
			738 => std_logic_vector(to_unsigned(247, 8)),
			739 => std_logic_vector(to_unsigned(30, 8)),
			740 => std_logic_vector(to_unsigned(128, 8)),
			741 => std_logic_vector(to_unsigned(208, 8)),
			742 => std_logic_vector(to_unsigned(68, 8)),
			743 => std_logic_vector(to_unsigned(183, 8)),
			744 => std_logic_vector(to_unsigned(183, 8)),
			745 => std_logic_vector(to_unsigned(169, 8)),
			746 => std_logic_vector(to_unsigned(75, 8)),
			747 => std_logic_vector(to_unsigned(186, 8)),
			748 => std_logic_vector(to_unsigned(31, 8)),
			749 => std_logic_vector(to_unsigned(126, 8)),
			750 => std_logic_vector(to_unsigned(217, 8)),
			751 => std_logic_vector(to_unsigned(31, 8)),
			752 => std_logic_vector(to_unsigned(61, 8)),
			753 => std_logic_vector(to_unsigned(134, 8)),
			754 => std_logic_vector(to_unsigned(177, 8)),
			755 => std_logic_vector(to_unsigned(189, 8)),
			756 => std_logic_vector(to_unsigned(192, 8)),
			757 => std_logic_vector(to_unsigned(145, 8)),
			758 => std_logic_vector(to_unsigned(156, 8)),
			759 => std_logic_vector(to_unsigned(72, 8)),
			760 => std_logic_vector(to_unsigned(211, 8)),
			761 => std_logic_vector(to_unsigned(116, 8)),
			762 => std_logic_vector(to_unsigned(234, 8)),
			763 => std_logic_vector(to_unsigned(210, 8)),
			764 => std_logic_vector(to_unsigned(234, 8)),
			765 => std_logic_vector(to_unsigned(175, 8)),
			766 => std_logic_vector(to_unsigned(186, 8)),
			767 => std_logic_vector(to_unsigned(208, 8)),
			768 => std_logic_vector(to_unsigned(22, 8)),
			769 => std_logic_vector(to_unsigned(33, 8)),
			770 => std_logic_vector(to_unsigned(7, 8)),
			771 => std_logic_vector(to_unsigned(250, 8)),
			772 => std_logic_vector(to_unsigned(196, 8)),
			773 => std_logic_vector(to_unsigned(168, 8)),
			774 => std_logic_vector(to_unsigned(102, 8)),
			775 => std_logic_vector(to_unsigned(88, 8)),
			776 => std_logic_vector(to_unsigned(106, 8)),
			777 => std_logic_vector(to_unsigned(57, 8)),
			778 => std_logic_vector(to_unsigned(0, 8)),
			779 => std_logic_vector(to_unsigned(95, 8)),
			780 => std_logic_vector(to_unsigned(127, 8)),
			781 => std_logic_vector(to_unsigned(177, 8)),
			782 => std_logic_vector(to_unsigned(138, 8)),
			783 => std_logic_vector(to_unsigned(165, 8)),
			784 => std_logic_vector(to_unsigned(187, 8)),
			785 => std_logic_vector(to_unsigned(19, 8)),
			786 => std_logic_vector(to_unsigned(221, 8)),
			787 => std_logic_vector(to_unsigned(160, 8)),
			788 => std_logic_vector(to_unsigned(46, 8)),
			789 => std_logic_vector(to_unsigned(47, 8)),
			790 => std_logic_vector(to_unsigned(73, 8)),
			791 => std_logic_vector(to_unsigned(144, 8)),
			792 => std_logic_vector(to_unsigned(131, 8)),
			793 => std_logic_vector(to_unsigned(2, 8)),
			794 => std_logic_vector(to_unsigned(124, 8)),
			795 => std_logic_vector(to_unsigned(16, 8)),
			796 => std_logic_vector(to_unsigned(220, 8)),
			797 => std_logic_vector(to_unsigned(214, 8)),
			798 => std_logic_vector(to_unsigned(143, 8)),
			799 => std_logic_vector(to_unsigned(188, 8)),
			800 => std_logic_vector(to_unsigned(131, 8)),
			801 => std_logic_vector(to_unsigned(239, 8)),
			802 => std_logic_vector(to_unsigned(201, 8)),
			803 => std_logic_vector(to_unsigned(44, 8)),
			804 => std_logic_vector(to_unsigned(137, 8)),
			805 => std_logic_vector(to_unsigned(155, 8)),
			806 => std_logic_vector(to_unsigned(220, 8)),
			807 => std_logic_vector(to_unsigned(232, 8)),
			808 => std_logic_vector(to_unsigned(82, 8)),
			809 => std_logic_vector(to_unsigned(114, 8)),
			810 => std_logic_vector(to_unsigned(80, 8)),
			811 => std_logic_vector(to_unsigned(24, 8)),
			812 => std_logic_vector(to_unsigned(102, 8)),
			813 => std_logic_vector(to_unsigned(93, 8)),
			814 => std_logic_vector(to_unsigned(0, 8)),
			815 => std_logic_vector(to_unsigned(59, 8)),
			816 => std_logic_vector(to_unsigned(55, 8)),
			817 => std_logic_vector(to_unsigned(118, 8)),
			818 => std_logic_vector(to_unsigned(7, 8)),
			819 => std_logic_vector(to_unsigned(139, 8)),
			820 => std_logic_vector(to_unsigned(222, 8)),
			821 => std_logic_vector(to_unsigned(224, 8)),
			822 => std_logic_vector(to_unsigned(236, 8)),
			823 => std_logic_vector(to_unsigned(75, 8)),
			824 => std_logic_vector(to_unsigned(92, 8)),
			825 => std_logic_vector(to_unsigned(199, 8)),
			826 => std_logic_vector(to_unsigned(119, 8)),
			827 => std_logic_vector(to_unsigned(56, 8)),
			828 => std_logic_vector(to_unsigned(224, 8)),
			829 => std_logic_vector(to_unsigned(42, 8)),
			830 => std_logic_vector(to_unsigned(152, 8)),
			831 => std_logic_vector(to_unsigned(249, 8)),
			832 => std_logic_vector(to_unsigned(25, 8)),
			833 => std_logic_vector(to_unsigned(197, 8)),
			834 => std_logic_vector(to_unsigned(247, 8)),
			835 => std_logic_vector(to_unsigned(152, 8)),
			836 => std_logic_vector(to_unsigned(60, 8)),
			837 => std_logic_vector(to_unsigned(107, 8)),
			838 => std_logic_vector(to_unsigned(183, 8)),
			839 => std_logic_vector(to_unsigned(185, 8)),
			840 => std_logic_vector(to_unsigned(79, 8)),
			841 => std_logic_vector(to_unsigned(231, 8)),
			842 => std_logic_vector(to_unsigned(149, 8)),
			843 => std_logic_vector(to_unsigned(31, 8)),
			844 => std_logic_vector(to_unsigned(31, 8)),
			845 => std_logic_vector(to_unsigned(215, 8)),
			846 => std_logic_vector(to_unsigned(25, 8)),
			847 => std_logic_vector(to_unsigned(4, 8)),
			848 => std_logic_vector(to_unsigned(58, 8)),
			849 => std_logic_vector(to_unsigned(8, 8)),
			850 => std_logic_vector(to_unsigned(188, 8)),
			851 => std_logic_vector(to_unsigned(56, 8)),
			852 => std_logic_vector(to_unsigned(188, 8)),
			853 => std_logic_vector(to_unsigned(1, 8)),
			854 => std_logic_vector(to_unsigned(17, 8)),
			855 => std_logic_vector(to_unsigned(9, 8)),
			856 => std_logic_vector(to_unsigned(203, 8)),
			857 => std_logic_vector(to_unsigned(192, 8)),
			858 => std_logic_vector(to_unsigned(12, 8)),
			859 => std_logic_vector(to_unsigned(70, 8)),
			860 => std_logic_vector(to_unsigned(12, 8)),
			861 => std_logic_vector(to_unsigned(133, 8)),
			862 => std_logic_vector(to_unsigned(156, 8)),
			863 => std_logic_vector(to_unsigned(207, 8)),
			864 => std_logic_vector(to_unsigned(46, 8)),
			865 => std_logic_vector(to_unsigned(70, 8)),
			866 => std_logic_vector(to_unsigned(89, 8)),
			867 => std_logic_vector(to_unsigned(93, 8)),
			868 => std_logic_vector(to_unsigned(255, 8)),
			869 => std_logic_vector(to_unsigned(226, 8)),
			870 => std_logic_vector(to_unsigned(32, 8)),
			871 => std_logic_vector(to_unsigned(34, 8)),
			872 => std_logic_vector(to_unsigned(192, 8)),
			873 => std_logic_vector(to_unsigned(33, 8)),
			874 => std_logic_vector(to_unsigned(154, 8)),
			875 => std_logic_vector(to_unsigned(27, 8)),
			876 => std_logic_vector(to_unsigned(90, 8)),
			877 => std_logic_vector(to_unsigned(248, 8)),
			878 => std_logic_vector(to_unsigned(175, 8)),
			879 => std_logic_vector(to_unsigned(49, 8)),
			880 => std_logic_vector(to_unsigned(82, 8)),
			881 => std_logic_vector(to_unsigned(219, 8)),
			882 => std_logic_vector(to_unsigned(67, 8)),
			883 => std_logic_vector(to_unsigned(9, 8)),
			884 => std_logic_vector(to_unsigned(229, 8)),
			885 => std_logic_vector(to_unsigned(125, 8)),
			886 => std_logic_vector(to_unsigned(196, 8)),
			887 => std_logic_vector(to_unsigned(196, 8)),
			888 => std_logic_vector(to_unsigned(102, 8)),
			889 => std_logic_vector(to_unsigned(165, 8)),
			890 => std_logic_vector(to_unsigned(209, 8)),
			891 => std_logic_vector(to_unsigned(152, 8)),
			892 => std_logic_vector(to_unsigned(117, 8)),
			893 => std_logic_vector(to_unsigned(174, 8)),
			894 => std_logic_vector(to_unsigned(117, 8)),
			895 => std_logic_vector(to_unsigned(164, 8)),
			896 => std_logic_vector(to_unsigned(9, 8)),
			897 => std_logic_vector(to_unsigned(108, 8)),
			898 => std_logic_vector(to_unsigned(154, 8)),
			899 => std_logic_vector(to_unsigned(76, 8)),
			900 => std_logic_vector(to_unsigned(210, 8)),
			901 => std_logic_vector(to_unsigned(149, 8)),
			902 => std_logic_vector(to_unsigned(230, 8)),
			903 => std_logic_vector(to_unsigned(79, 8)),
			904 => std_logic_vector(to_unsigned(95, 8)),
			905 => std_logic_vector(to_unsigned(81, 8)),
			906 => std_logic_vector(to_unsigned(2, 8)),
			907 => std_logic_vector(to_unsigned(138, 8)),
			908 => std_logic_vector(to_unsigned(8, 8)),
			909 => std_logic_vector(to_unsigned(195, 8)),
			910 => std_logic_vector(to_unsigned(65, 8)),
			911 => std_logic_vector(to_unsigned(245, 8)),
			912 => std_logic_vector(to_unsigned(206, 8)),
			913 => std_logic_vector(to_unsigned(2, 8)),
			914 => std_logic_vector(to_unsigned(187, 8)),
			915 => std_logic_vector(to_unsigned(192, 8)),
			916 => std_logic_vector(to_unsigned(242, 8)),
			917 => std_logic_vector(to_unsigned(52, 8)),
			918 => std_logic_vector(to_unsigned(81, 8)),
			919 => std_logic_vector(to_unsigned(110, 8)),
			920 => std_logic_vector(to_unsigned(105, 8)),
			921 => std_logic_vector(to_unsigned(1, 8)),
			922 => std_logic_vector(to_unsigned(214, 8)),
			923 => std_logic_vector(to_unsigned(2, 8)),
			924 => std_logic_vector(to_unsigned(246, 8)),
			925 => std_logic_vector(to_unsigned(248, 8)),
			926 => std_logic_vector(to_unsigned(106, 8)),
			927 => std_logic_vector(to_unsigned(138, 8)),
			928 => std_logic_vector(to_unsigned(47, 8)),
			929 => std_logic_vector(to_unsigned(211, 8)),
			930 => std_logic_vector(to_unsigned(139, 8)),
			931 => std_logic_vector(to_unsigned(180, 8)),
			932 => std_logic_vector(to_unsigned(2, 8)),
			933 => std_logic_vector(to_unsigned(78, 8)),
			934 => std_logic_vector(to_unsigned(42, 8)),
			935 => std_logic_vector(to_unsigned(92, 8)),
			936 => std_logic_vector(to_unsigned(43, 8)),
			937 => std_logic_vector(to_unsigned(157, 8)),
			938 => std_logic_vector(to_unsigned(80, 8)),
			939 => std_logic_vector(to_unsigned(97, 8)),
			940 => std_logic_vector(to_unsigned(216, 8)),
			941 => std_logic_vector(to_unsigned(14, 8)),
			942 => std_logic_vector(to_unsigned(43, 8)),
			943 => std_logic_vector(to_unsigned(247, 8)),
			944 => std_logic_vector(to_unsigned(140, 8)),
			945 => std_logic_vector(to_unsigned(102, 8)),
			946 => std_logic_vector(to_unsigned(151, 8)),
			947 => std_logic_vector(to_unsigned(137, 8)),
			948 => std_logic_vector(to_unsigned(102, 8)),
			949 => std_logic_vector(to_unsigned(39, 8)),
			950 => std_logic_vector(to_unsigned(66, 8)),
			951 => std_logic_vector(to_unsigned(102, 8)),
			952 => std_logic_vector(to_unsigned(146, 8)),
			953 => std_logic_vector(to_unsigned(211, 8)),
			954 => std_logic_vector(to_unsigned(108, 8)),
			955 => std_logic_vector(to_unsigned(104, 8)),
			956 => std_logic_vector(to_unsigned(22, 8)),
			957 => std_logic_vector(to_unsigned(86, 8)),
			958 => std_logic_vector(to_unsigned(112, 8)),
			959 => std_logic_vector(to_unsigned(9, 8)),
			960 => std_logic_vector(to_unsigned(112, 8)),
			961 => std_logic_vector(to_unsigned(48, 8)),
			962 => std_logic_vector(to_unsigned(29, 8)),
			963 => std_logic_vector(to_unsigned(32, 8)),
			964 => std_logic_vector(to_unsigned(154, 8)),
			965 => std_logic_vector(to_unsigned(76, 8)),
			966 => std_logic_vector(to_unsigned(69, 8)),
			967 => std_logic_vector(to_unsigned(37, 8)),
			968 => std_logic_vector(to_unsigned(41, 8)),
			969 => std_logic_vector(to_unsigned(122, 8)),
			970 => std_logic_vector(to_unsigned(74, 8)),
			971 => std_logic_vector(to_unsigned(137, 8)),
			972 => std_logic_vector(to_unsigned(154, 8)),
			973 => std_logic_vector(to_unsigned(185, 8)),
			974 => std_logic_vector(to_unsigned(173, 8)),
			975 => std_logic_vector(to_unsigned(18, 8)),
			976 => std_logic_vector(to_unsigned(169, 8)),
			977 => std_logic_vector(to_unsigned(77, 8)),
			978 => std_logic_vector(to_unsigned(208, 8)),
			979 => std_logic_vector(to_unsigned(65, 8)),
			980 => std_logic_vector(to_unsigned(25, 8)),
			981 => std_logic_vector(to_unsigned(251, 8)),
			982 => std_logic_vector(to_unsigned(73, 8)),
			983 => std_logic_vector(to_unsigned(168, 8)),
			984 => std_logic_vector(to_unsigned(125, 8)),
			985 => std_logic_vector(to_unsigned(63, 8)),
			986 => std_logic_vector(to_unsigned(93, 8)),
			987 => std_logic_vector(to_unsigned(235, 8)),
			988 => std_logic_vector(to_unsigned(253, 8)),
			989 => std_logic_vector(to_unsigned(24, 8)),
			990 => std_logic_vector(to_unsigned(10, 8)),
			991 => std_logic_vector(to_unsigned(133, 8)),
			992 => std_logic_vector(to_unsigned(178, 8)),
			993 => std_logic_vector(to_unsigned(237, 8)),
			994 => std_logic_vector(to_unsigned(72, 8)),
			995 => std_logic_vector(to_unsigned(178, 8)),
			996 => std_logic_vector(to_unsigned(183, 8)),
			997 => std_logic_vector(to_unsigned(203, 8)),
			998 => std_logic_vector(to_unsigned(21, 8)),
			999 => std_logic_vector(to_unsigned(254, 8)),
			1000 => std_logic_vector(to_unsigned(87, 8)),
			1001 => std_logic_vector(to_unsigned(82, 8)),
			1002 => std_logic_vector(to_unsigned(76, 8)),
			1003 => std_logic_vector(to_unsigned(192, 8)),
			1004 => std_logic_vector(to_unsigned(14, 8)),
			1005 => std_logic_vector(to_unsigned(108, 8)),
			1006 => std_logic_vector(to_unsigned(218, 8)),
			1007 => std_logic_vector(to_unsigned(196, 8)),
			1008 => std_logic_vector(to_unsigned(8, 8)),
			1009 => std_logic_vector(to_unsigned(4, 8)),
			1010 => std_logic_vector(to_unsigned(224, 8)),
			1011 => std_logic_vector(to_unsigned(48, 8)),
			1012 => std_logic_vector(to_unsigned(93, 8)),
			1013 => std_logic_vector(to_unsigned(64, 8)),
			1014 => std_logic_vector(to_unsigned(228, 8)),
			1015 => std_logic_vector(to_unsigned(206, 8)),
			1016 => std_logic_vector(to_unsigned(225, 8)),
			1017 => std_logic_vector(to_unsigned(189, 8)),
			1018 => std_logic_vector(to_unsigned(126, 8)),
			1019 => std_logic_vector(to_unsigned(47, 8)),
			1020 => std_logic_vector(to_unsigned(173, 8)),
			1021 => std_logic_vector(to_unsigned(243, 8)),
			1022 => std_logic_vector(to_unsigned(5, 8)),
			1023 => std_logic_vector(to_unsigned(75, 8)),
			1024 => std_logic_vector(to_unsigned(163, 8)),
			1025 => std_logic_vector(to_unsigned(132, 8)),
			1026 => std_logic_vector(to_unsigned(231, 8)),
			1027 => std_logic_vector(to_unsigned(33, 8)),
			1028 => std_logic_vector(to_unsigned(23, 8)),
			1029 => std_logic_vector(to_unsigned(111, 8)),
			1030 => std_logic_vector(to_unsigned(85, 8)),
			1031 => std_logic_vector(to_unsigned(121, 8)),
			1032 => std_logic_vector(to_unsigned(171, 8)),
			1033 => std_logic_vector(to_unsigned(79, 8)),
			1034 => std_logic_vector(to_unsigned(111, 8)),
			1035 => std_logic_vector(to_unsigned(220, 8)),
			1036 => std_logic_vector(to_unsigned(249, 8)),
			1037 => std_logic_vector(to_unsigned(241, 8)),
			1038 => std_logic_vector(to_unsigned(219, 8)),
			1039 => std_logic_vector(to_unsigned(16, 8)),
			1040 => std_logic_vector(to_unsigned(212, 8)),
			1041 => std_logic_vector(to_unsigned(7, 8)),
			1042 => std_logic_vector(to_unsigned(92, 8)),
			1043 => std_logic_vector(to_unsigned(15, 8)),
			1044 => std_logic_vector(to_unsigned(125, 8)),
			1045 => std_logic_vector(to_unsigned(89, 8)),
			1046 => std_logic_vector(to_unsigned(39, 8)),
			1047 => std_logic_vector(to_unsigned(68, 8)),
			1048 => std_logic_vector(to_unsigned(27, 8)),
			1049 => std_logic_vector(to_unsigned(178, 8)),
			1050 => std_logic_vector(to_unsigned(213, 8)),
			1051 => std_logic_vector(to_unsigned(212, 8)),
			1052 => std_logic_vector(to_unsigned(235, 8)),
			1053 => std_logic_vector(to_unsigned(10, 8)),
			1054 => std_logic_vector(to_unsigned(173, 8)),
			1055 => std_logic_vector(to_unsigned(79, 8)),
			1056 => std_logic_vector(to_unsigned(226, 8)),
			1057 => std_logic_vector(to_unsigned(197, 8)),
			1058 => std_logic_vector(to_unsigned(240, 8)),
			1059 => std_logic_vector(to_unsigned(175, 8)),
			1060 => std_logic_vector(to_unsigned(69, 8)),
			1061 => std_logic_vector(to_unsigned(183, 8)),
			1062 => std_logic_vector(to_unsigned(121, 8)),
			1063 => std_logic_vector(to_unsigned(189, 8)),
			1064 => std_logic_vector(to_unsigned(171, 8)),
			1065 => std_logic_vector(to_unsigned(101, 8)),
			1066 => std_logic_vector(to_unsigned(6, 8)),
			1067 => std_logic_vector(to_unsigned(100, 8)),
			1068 => std_logic_vector(to_unsigned(247, 8)),
			1069 => std_logic_vector(to_unsigned(91, 8)),
			1070 => std_logic_vector(to_unsigned(233, 8)),
			1071 => std_logic_vector(to_unsigned(227, 8)),
			1072 => std_logic_vector(to_unsigned(76, 8)),
			1073 => std_logic_vector(to_unsigned(106, 8)),
			1074 => std_logic_vector(to_unsigned(184, 8)),
			1075 => std_logic_vector(to_unsigned(76, 8)),
			1076 => std_logic_vector(to_unsigned(4, 8)),
			1077 => std_logic_vector(to_unsigned(110, 8)),
			1078 => std_logic_vector(to_unsigned(41, 8)),
			1079 => std_logic_vector(to_unsigned(214, 8)),
			1080 => std_logic_vector(to_unsigned(86, 8)),
			1081 => std_logic_vector(to_unsigned(112, 8)),
			1082 => std_logic_vector(to_unsigned(34, 8)),
			1083 => std_logic_vector(to_unsigned(162, 8)),
			1084 => std_logic_vector(to_unsigned(31, 8)),
			1085 => std_logic_vector(to_unsigned(0, 8)),
			1086 => std_logic_vector(to_unsigned(65, 8)),
			1087 => std_logic_vector(to_unsigned(171, 8)),
			1088 => std_logic_vector(to_unsigned(227, 8)),
			1089 => std_logic_vector(to_unsigned(166, 8)),
			1090 => std_logic_vector(to_unsigned(245, 8)),
			1091 => std_logic_vector(to_unsigned(160, 8)),
			1092 => std_logic_vector(to_unsigned(56, 8)),
			1093 => std_logic_vector(to_unsigned(241, 8)),
			1094 => std_logic_vector(to_unsigned(241, 8)),
			1095 => std_logic_vector(to_unsigned(97, 8)),
			1096 => std_logic_vector(to_unsigned(95, 8)),
			1097 => std_logic_vector(to_unsigned(31, 8)),
			1098 => std_logic_vector(to_unsigned(59, 8)),
			1099 => std_logic_vector(to_unsigned(137, 8)),
			1100 => std_logic_vector(to_unsigned(134, 8)),
			1101 => std_logic_vector(to_unsigned(166, 8)),
			1102 => std_logic_vector(to_unsigned(227, 8)),
			1103 => std_logic_vector(to_unsigned(213, 8)),
			1104 => std_logic_vector(to_unsigned(92, 8)),
			1105 => std_logic_vector(to_unsigned(14, 8)),
			1106 => std_logic_vector(to_unsigned(68, 8)),
			1107 => std_logic_vector(to_unsigned(115, 8)),
			1108 => std_logic_vector(to_unsigned(82, 8)),
			1109 => std_logic_vector(to_unsigned(165, 8)),
			1110 => std_logic_vector(to_unsigned(252, 8)),
			1111 => std_logic_vector(to_unsigned(187, 8)),
			1112 => std_logic_vector(to_unsigned(60, 8)),
			1113 => std_logic_vector(to_unsigned(170, 8)),
			1114 => std_logic_vector(to_unsigned(242, 8)),
			1115 => std_logic_vector(to_unsigned(174, 8)),
			1116 => std_logic_vector(to_unsigned(93, 8)),
			1117 => std_logic_vector(to_unsigned(15, 8)),
			1118 => std_logic_vector(to_unsigned(213, 8)),
			1119 => std_logic_vector(to_unsigned(28, 8)),
			1120 => std_logic_vector(to_unsigned(45, 8)),
			1121 => std_logic_vector(to_unsigned(15, 8)),
			1122 => std_logic_vector(to_unsigned(226, 8)),
			1123 => std_logic_vector(to_unsigned(208, 8)),
			1124 => std_logic_vector(to_unsigned(87, 8)),
			1125 => std_logic_vector(to_unsigned(126, 8)),
			1126 => std_logic_vector(to_unsigned(38, 8)),
			1127 => std_logic_vector(to_unsigned(7, 8)),
			1128 => std_logic_vector(to_unsigned(173, 8)),
			1129 => std_logic_vector(to_unsigned(206, 8)),
			1130 => std_logic_vector(to_unsigned(110, 8)),
			1131 => std_logic_vector(to_unsigned(204, 8)),
			1132 => std_logic_vector(to_unsigned(34, 8)),
			1133 => std_logic_vector(to_unsigned(233, 8)),
			1134 => std_logic_vector(to_unsigned(234, 8)),
			1135 => std_logic_vector(to_unsigned(213, 8)),
			1136 => std_logic_vector(to_unsigned(139, 8)),
			1137 => std_logic_vector(to_unsigned(221, 8)),
			1138 => std_logic_vector(to_unsigned(86, 8)),
			1139 => std_logic_vector(to_unsigned(218, 8)),
			1140 => std_logic_vector(to_unsigned(3, 8)),
			1141 => std_logic_vector(to_unsigned(48, 8)),
			1142 => std_logic_vector(to_unsigned(21, 8)),
			1143 => std_logic_vector(to_unsigned(239, 8)),
			1144 => std_logic_vector(to_unsigned(131, 8)),
			1145 => std_logic_vector(to_unsigned(190, 8)),
			1146 => std_logic_vector(to_unsigned(80, 8)),
			1147 => std_logic_vector(to_unsigned(108, 8)),
			1148 => std_logic_vector(to_unsigned(188, 8)),
			1149 => std_logic_vector(to_unsigned(151, 8)),
			1150 => std_logic_vector(to_unsigned(215, 8)),
			1151 => std_logic_vector(to_unsigned(21, 8)),
			1152 => std_logic_vector(to_unsigned(245, 8)),
			1153 => std_logic_vector(to_unsigned(36, 8)),
			1154 => std_logic_vector(to_unsigned(182, 8)),
			1155 => std_logic_vector(to_unsigned(143, 8)),
			1156 => std_logic_vector(to_unsigned(245, 8)),
			1157 => std_logic_vector(to_unsigned(189, 8)),
			1158 => std_logic_vector(to_unsigned(149, 8)),
			1159 => std_logic_vector(to_unsigned(158, 8)),
			1160 => std_logic_vector(to_unsigned(251, 8)),
			1161 => std_logic_vector(to_unsigned(248, 8)),
			1162 => std_logic_vector(to_unsigned(147, 8)),
			1163 => std_logic_vector(to_unsigned(140, 8)),
			1164 => std_logic_vector(to_unsigned(178, 8)),
			1165 => std_logic_vector(to_unsigned(167, 8)),
			1166 => std_logic_vector(to_unsigned(144, 8)),
			1167 => std_logic_vector(to_unsigned(78, 8)),
			1168 => std_logic_vector(to_unsigned(63, 8)),
			1169 => std_logic_vector(to_unsigned(213, 8)),
			1170 => std_logic_vector(to_unsigned(83, 8)),
			1171 => std_logic_vector(to_unsigned(163, 8)),
			1172 => std_logic_vector(to_unsigned(10, 8)),
			1173 => std_logic_vector(to_unsigned(212, 8)),
			1174 => std_logic_vector(to_unsigned(188, 8)),
			1175 => std_logic_vector(to_unsigned(104, 8)),
			1176 => std_logic_vector(to_unsigned(187, 8)),
			1177 => std_logic_vector(to_unsigned(153, 8)),
			1178 => std_logic_vector(to_unsigned(32, 8)),
			1179 => std_logic_vector(to_unsigned(112, 8)),
			1180 => std_logic_vector(to_unsigned(88, 8)),
			1181 => std_logic_vector(to_unsigned(176, 8)),
			1182 => std_logic_vector(to_unsigned(135, 8)),
			1183 => std_logic_vector(to_unsigned(10, 8)),
			1184 => std_logic_vector(to_unsigned(108, 8)),
			1185 => std_logic_vector(to_unsigned(201, 8)),
			1186 => std_logic_vector(to_unsigned(182, 8)),
			1187 => std_logic_vector(to_unsigned(140, 8)),
			1188 => std_logic_vector(to_unsigned(10, 8)),
			1189 => std_logic_vector(to_unsigned(144, 8)),
			1190 => std_logic_vector(to_unsigned(49, 8)),
			1191 => std_logic_vector(to_unsigned(124, 8)),
			1192 => std_logic_vector(to_unsigned(207, 8)),
			1193 => std_logic_vector(to_unsigned(7, 8)),
			1194 => std_logic_vector(to_unsigned(229, 8)),
			1195 => std_logic_vector(to_unsigned(44, 8)),
			1196 => std_logic_vector(to_unsigned(193, 8)),
			1197 => std_logic_vector(to_unsigned(22, 8)),
			1198 => std_logic_vector(to_unsigned(240, 8)),
			1199 => std_logic_vector(to_unsigned(85, 8)),
			1200 => std_logic_vector(to_unsigned(109, 8)),
			1201 => std_logic_vector(to_unsigned(194, 8)),
			1202 => std_logic_vector(to_unsigned(202, 8)),
			1203 => std_logic_vector(to_unsigned(117, 8)),
			1204 => std_logic_vector(to_unsigned(201, 8)),
			1205 => std_logic_vector(to_unsigned(122, 8)),
			1206 => std_logic_vector(to_unsigned(194, 8)),
			1207 => std_logic_vector(to_unsigned(81, 8)),
			1208 => std_logic_vector(to_unsigned(15, 8)),
			1209 => std_logic_vector(to_unsigned(154, 8)),
			1210 => std_logic_vector(to_unsigned(162, 8)),
			1211 => std_logic_vector(to_unsigned(36, 8)),
			1212 => std_logic_vector(to_unsigned(213, 8)),
			1213 => std_logic_vector(to_unsigned(187, 8)),
			1214 => std_logic_vector(to_unsigned(202, 8)),
			1215 => std_logic_vector(to_unsigned(108, 8)),
			1216 => std_logic_vector(to_unsigned(232, 8)),
			1217 => std_logic_vector(to_unsigned(137, 8)),
			1218 => std_logic_vector(to_unsigned(232, 8)),
			1219 => std_logic_vector(to_unsigned(189, 8)),
			1220 => std_logic_vector(to_unsigned(218, 8)),
			1221 => std_logic_vector(to_unsigned(66, 8)),
			1222 => std_logic_vector(to_unsigned(168, 8)),
			1223 => std_logic_vector(to_unsigned(144, 8)),
			1224 => std_logic_vector(to_unsigned(71, 8)),
			1225 => std_logic_vector(to_unsigned(120, 8)),
			1226 => std_logic_vector(to_unsigned(240, 8)),
			1227 => std_logic_vector(to_unsigned(91, 8)),
			1228 => std_logic_vector(to_unsigned(32, 8)),
			1229 => std_logic_vector(to_unsigned(84, 8)),
			1230 => std_logic_vector(to_unsigned(173, 8)),
			1231 => std_logic_vector(to_unsigned(189, 8)),
			1232 => std_logic_vector(to_unsigned(67, 8)),
			1233 => std_logic_vector(to_unsigned(196, 8)),
			1234 => std_logic_vector(to_unsigned(27, 8)),
			1235 => std_logic_vector(to_unsigned(18, 8)),
			1236 => std_logic_vector(to_unsigned(183, 8)),
			1237 => std_logic_vector(to_unsigned(79, 8)),
			1238 => std_logic_vector(to_unsigned(22, 8)),
			1239 => std_logic_vector(to_unsigned(125, 8)),
			1240 => std_logic_vector(to_unsigned(32, 8)),
			1241 => std_logic_vector(to_unsigned(98, 8)),
			1242 => std_logic_vector(to_unsigned(39, 8)),
			1243 => std_logic_vector(to_unsigned(67, 8)),
			1244 => std_logic_vector(to_unsigned(116, 8)),
			1245 => std_logic_vector(to_unsigned(43, 8)),
			1246 => std_logic_vector(to_unsigned(103, 8)),
			1247 => std_logic_vector(to_unsigned(226, 8)),
			1248 => std_logic_vector(to_unsigned(10, 8)),
			1249 => std_logic_vector(to_unsigned(225, 8)),
			1250 => std_logic_vector(to_unsigned(98, 8)),
			1251 => std_logic_vector(to_unsigned(29, 8)),
			1252 => std_logic_vector(to_unsigned(225, 8)),
			1253 => std_logic_vector(to_unsigned(39, 8)),
			1254 => std_logic_vector(to_unsigned(152, 8)),
			1255 => std_logic_vector(to_unsigned(187, 8)),
			1256 => std_logic_vector(to_unsigned(93, 8)),
			1257 => std_logic_vector(to_unsigned(27, 8)),
			1258 => std_logic_vector(to_unsigned(26, 8)),
			1259 => std_logic_vector(to_unsigned(39, 8)),
			1260 => std_logic_vector(to_unsigned(17, 8)),
			1261 => std_logic_vector(to_unsigned(38, 8)),
			1262 => std_logic_vector(to_unsigned(117, 8)),
			1263 => std_logic_vector(to_unsigned(85, 8)),
			1264 => std_logic_vector(to_unsigned(117, 8)),
			1265 => std_logic_vector(to_unsigned(115, 8)),
			1266 => std_logic_vector(to_unsigned(11, 8)),
			1267 => std_logic_vector(to_unsigned(148, 8)),
			1268 => std_logic_vector(to_unsigned(167, 8)),
			1269 => std_logic_vector(to_unsigned(117, 8)),
			1270 => std_logic_vector(to_unsigned(11, 8)),
			1271 => std_logic_vector(to_unsigned(208, 8)),
			1272 => std_logic_vector(to_unsigned(78, 8)),
			1273 => std_logic_vector(to_unsigned(103, 8)),
			1274 => std_logic_vector(to_unsigned(40, 8)),
			1275 => std_logic_vector(to_unsigned(92, 8)),
			1276 => std_logic_vector(to_unsigned(6, 8)),
			1277 => std_logic_vector(to_unsigned(62, 8)),
			1278 => std_logic_vector(to_unsigned(30, 8)),
			1279 => std_logic_vector(to_unsigned(143, 8)),
			1280 => std_logic_vector(to_unsigned(65, 8)),
			1281 => std_logic_vector(to_unsigned(137, 8)),
			1282 => std_logic_vector(to_unsigned(48, 8)),
			1283 => std_logic_vector(to_unsigned(179, 8)),
			1284 => std_logic_vector(to_unsigned(51, 8)),
			1285 => std_logic_vector(to_unsigned(247, 8)),
			1286 => std_logic_vector(to_unsigned(104, 8)),
			1287 => std_logic_vector(to_unsigned(98, 8)),
			1288 => std_logic_vector(to_unsigned(181, 8)),
			1289 => std_logic_vector(to_unsigned(12, 8)),
			1290 => std_logic_vector(to_unsigned(85, 8)),
			1291 => std_logic_vector(to_unsigned(173, 8)),
			1292 => std_logic_vector(to_unsigned(216, 8)),
			1293 => std_logic_vector(to_unsigned(71, 8)),
			1294 => std_logic_vector(to_unsigned(116, 8)),
			1295 => std_logic_vector(to_unsigned(197, 8)),
			1296 => std_logic_vector(to_unsigned(167, 8)),
			1297 => std_logic_vector(to_unsigned(156, 8)),
			1298 => std_logic_vector(to_unsigned(4, 8)),
			1299 => std_logic_vector(to_unsigned(86, 8)),
			1300 => std_logic_vector(to_unsigned(77, 8)),
			1301 => std_logic_vector(to_unsigned(169, 8)),
			1302 => std_logic_vector(to_unsigned(58, 8)),
			1303 => std_logic_vector(to_unsigned(174, 8)),
			1304 => std_logic_vector(to_unsigned(139, 8)),
			1305 => std_logic_vector(to_unsigned(117, 8)),
			1306 => std_logic_vector(to_unsigned(131, 8)),
			1307 => std_logic_vector(to_unsigned(86, 8)),
			1308 => std_logic_vector(to_unsigned(162, 8)),
			1309 => std_logic_vector(to_unsigned(79, 8)),
			1310 => std_logic_vector(to_unsigned(153, 8)),
			1311 => std_logic_vector(to_unsigned(156, 8)),
			1312 => std_logic_vector(to_unsigned(212, 8)),
			1313 => std_logic_vector(to_unsigned(248, 8)),
			1314 => std_logic_vector(to_unsigned(1, 8)),
			1315 => std_logic_vector(to_unsigned(12, 8)),
			1316 => std_logic_vector(to_unsigned(146, 8)),
			1317 => std_logic_vector(to_unsigned(191, 8)),
			1318 => std_logic_vector(to_unsigned(25, 8)),
			1319 => std_logic_vector(to_unsigned(19, 8)),
			1320 => std_logic_vector(to_unsigned(236, 8)),
			1321 => std_logic_vector(to_unsigned(26, 8)),
			1322 => std_logic_vector(to_unsigned(90, 8)),
			1323 => std_logic_vector(to_unsigned(2, 8)),
			1324 => std_logic_vector(to_unsigned(118, 8)),
			1325 => std_logic_vector(to_unsigned(33, 8)),
			1326 => std_logic_vector(to_unsigned(134, 8)),
			1327 => std_logic_vector(to_unsigned(1, 8)),
			1328 => std_logic_vector(to_unsigned(14, 8)),
			1329 => std_logic_vector(to_unsigned(156, 8)),
			1330 => std_logic_vector(to_unsigned(99, 8)),
			1331 => std_logic_vector(to_unsigned(176, 8)),
			1332 => std_logic_vector(to_unsigned(4, 8)),
			1333 => std_logic_vector(to_unsigned(34, 8)),
			1334 => std_logic_vector(to_unsigned(92, 8)),
			1335 => std_logic_vector(to_unsigned(67, 8)),
			1336 => std_logic_vector(to_unsigned(34, 8)),
			1337 => std_logic_vector(to_unsigned(254, 8)),
			1338 => std_logic_vector(to_unsigned(243, 8)),
			1339 => std_logic_vector(to_unsigned(58, 8)),
			1340 => std_logic_vector(to_unsigned(239, 8)),
			1341 => std_logic_vector(to_unsigned(112, 8)),
			1342 => std_logic_vector(to_unsigned(232, 8)),
			1343 => std_logic_vector(to_unsigned(154, 8)),
			1344 => std_logic_vector(to_unsigned(156, 8)),
			1345 => std_logic_vector(to_unsigned(47, 8)),
			1346 => std_logic_vector(to_unsigned(25, 8)),
			1347 => std_logic_vector(to_unsigned(83, 8)),
			1348 => std_logic_vector(to_unsigned(231, 8)),
			1349 => std_logic_vector(to_unsigned(225, 8)),
			1350 => std_logic_vector(to_unsigned(53, 8)),
			1351 => std_logic_vector(to_unsigned(8, 8)),
			1352 => std_logic_vector(to_unsigned(78, 8)),
			1353 => std_logic_vector(to_unsigned(148, 8)),
			1354 => std_logic_vector(to_unsigned(230, 8)),
			1355 => std_logic_vector(to_unsigned(86, 8)),
			1356 => std_logic_vector(to_unsigned(124, 8)),
			1357 => std_logic_vector(to_unsigned(170, 8)),
			1358 => std_logic_vector(to_unsigned(187, 8)),
			1359 => std_logic_vector(to_unsigned(24, 8)),
			1360 => std_logic_vector(to_unsigned(72, 8)),
			1361 => std_logic_vector(to_unsigned(7, 8)),
			1362 => std_logic_vector(to_unsigned(174, 8)),
			1363 => std_logic_vector(to_unsigned(161, 8)),
			1364 => std_logic_vector(to_unsigned(190, 8)),
			1365 => std_logic_vector(to_unsigned(96, 8)),
			1366 => std_logic_vector(to_unsigned(19, 8)),
			1367 => std_logic_vector(to_unsigned(217, 8)),
			1368 => std_logic_vector(to_unsigned(195, 8)),
			1369 => std_logic_vector(to_unsigned(45, 8)),
			1370 => std_logic_vector(to_unsigned(57, 8)),
			1371 => std_logic_vector(to_unsigned(151, 8)),
			1372 => std_logic_vector(to_unsigned(77, 8)),
			1373 => std_logic_vector(to_unsigned(203, 8)),
			1374 => std_logic_vector(to_unsigned(187, 8)),
			1375 => std_logic_vector(to_unsigned(36, 8)),
			1376 => std_logic_vector(to_unsigned(88, 8)),
			1377 => std_logic_vector(to_unsigned(160, 8)),
			1378 => std_logic_vector(to_unsigned(134, 8)),
			1379 => std_logic_vector(to_unsigned(95, 8)),
			1380 => std_logic_vector(to_unsigned(16, 8)),
			1381 => std_logic_vector(to_unsigned(230, 8)),
			1382 => std_logic_vector(to_unsigned(213, 8)),
			1383 => std_logic_vector(to_unsigned(129, 8)),
			1384 => std_logic_vector(to_unsigned(51, 8)),
			1385 => std_logic_vector(to_unsigned(176, 8)),
			1386 => std_logic_vector(to_unsigned(18, 8)),
			1387 => std_logic_vector(to_unsigned(248, 8)),
			1388 => std_logic_vector(to_unsigned(58, 8)),
			1389 => std_logic_vector(to_unsigned(167, 8)),
			1390 => std_logic_vector(to_unsigned(68, 8)),
			1391 => std_logic_vector(to_unsigned(92, 8)),
			1392 => std_logic_vector(to_unsigned(241, 8)),
			1393 => std_logic_vector(to_unsigned(84, 8)),
			1394 => std_logic_vector(to_unsigned(107, 8)),
			1395 => std_logic_vector(to_unsigned(245, 8)),
			1396 => std_logic_vector(to_unsigned(254, 8)),
			1397 => std_logic_vector(to_unsigned(169, 8)),
			1398 => std_logic_vector(to_unsigned(117, 8)),
			1399 => std_logic_vector(to_unsigned(136, 8)),
			1400 => std_logic_vector(to_unsigned(219, 8)),
			1401 => std_logic_vector(to_unsigned(244, 8)),
			1402 => std_logic_vector(to_unsigned(42, 8)),
			1403 => std_logic_vector(to_unsigned(160, 8)),
			1404 => std_logic_vector(to_unsigned(5, 8)),
			1405 => std_logic_vector(to_unsigned(8, 8)),
			1406 => std_logic_vector(to_unsigned(11, 8)),
			1407 => std_logic_vector(to_unsigned(103, 8)),
			1408 => std_logic_vector(to_unsigned(154, 8)),
			1409 => std_logic_vector(to_unsigned(174, 8)),
			1410 => std_logic_vector(to_unsigned(211, 8)),
			1411 => std_logic_vector(to_unsigned(115, 8)),
			1412 => std_logic_vector(to_unsigned(183, 8)),
			1413 => std_logic_vector(to_unsigned(1, 8)),
			1414 => std_logic_vector(to_unsigned(117, 8)),
			1415 => std_logic_vector(to_unsigned(18, 8)),
			1416 => std_logic_vector(to_unsigned(148, 8)),
			1417 => std_logic_vector(to_unsigned(38, 8)),
			1418 => std_logic_vector(to_unsigned(131, 8)),
			1419 => std_logic_vector(to_unsigned(40, 8)),
			1420 => std_logic_vector(to_unsigned(152, 8)),
			1421 => std_logic_vector(to_unsigned(229, 8)),
			1422 => std_logic_vector(to_unsigned(64, 8)),
			1423 => std_logic_vector(to_unsigned(80, 8)),
			1424 => std_logic_vector(to_unsigned(204, 8)),
			1425 => std_logic_vector(to_unsigned(61, 8)),
			1426 => std_logic_vector(to_unsigned(139, 8)),
			1427 => std_logic_vector(to_unsigned(78, 8)),
			1428 => std_logic_vector(to_unsigned(42, 8)),
			1429 => std_logic_vector(to_unsigned(78, 8)),
			1430 => std_logic_vector(to_unsigned(161, 8)),
			1431 => std_logic_vector(to_unsigned(253, 8)),
			1432 => std_logic_vector(to_unsigned(174, 8)),
			1433 => std_logic_vector(to_unsigned(59, 8)),
			1434 => std_logic_vector(to_unsigned(71, 8)),
			1435 => std_logic_vector(to_unsigned(44, 8)),
			1436 => std_logic_vector(to_unsigned(218, 8)),
			1437 => std_logic_vector(to_unsigned(158, 8)),
			1438 => std_logic_vector(to_unsigned(255, 8)),
			1439 => std_logic_vector(to_unsigned(214, 8)),
			1440 => std_logic_vector(to_unsigned(138, 8)),
			1441 => std_logic_vector(to_unsigned(176, 8)),
			1442 => std_logic_vector(to_unsigned(242, 8)),
			1443 => std_logic_vector(to_unsigned(239, 8)),
			1444 => std_logic_vector(to_unsigned(246, 8)),
			1445 => std_logic_vector(to_unsigned(157, 8)),
			1446 => std_logic_vector(to_unsigned(12, 8)),
			1447 => std_logic_vector(to_unsigned(22, 8)),
			1448 => std_logic_vector(to_unsigned(239, 8)),
			1449 => std_logic_vector(to_unsigned(163, 8)),
			1450 => std_logic_vector(to_unsigned(9, 8)),
			1451 => std_logic_vector(to_unsigned(246, 8)),
			1452 => std_logic_vector(to_unsigned(200, 8)),
			1453 => std_logic_vector(to_unsigned(45, 8)),
			1454 => std_logic_vector(to_unsigned(224, 8)),
			1455 => std_logic_vector(to_unsigned(20, 8)),
			1456 => std_logic_vector(to_unsigned(185, 8)),
			1457 => std_logic_vector(to_unsigned(87, 8)),
			1458 => std_logic_vector(to_unsigned(79, 8)),
			1459 => std_logic_vector(to_unsigned(38, 8)),
			1460 => std_logic_vector(to_unsigned(95, 8)),
			1461 => std_logic_vector(to_unsigned(137, 8)),
			1462 => std_logic_vector(to_unsigned(215, 8)),
			1463 => std_logic_vector(to_unsigned(252, 8)),
			1464 => std_logic_vector(to_unsigned(165, 8)),
			1465 => std_logic_vector(to_unsigned(16, 8)),
			1466 => std_logic_vector(to_unsigned(238, 8)),
			1467 => std_logic_vector(to_unsigned(137, 8)),
			1468 => std_logic_vector(to_unsigned(228, 8)),
			1469 => std_logic_vector(to_unsigned(75, 8)),
			1470 => std_logic_vector(to_unsigned(29, 8)),
			1471 => std_logic_vector(to_unsigned(97, 8)),
			1472 => std_logic_vector(to_unsigned(148, 8)),
			1473 => std_logic_vector(to_unsigned(112, 8)),
			1474 => std_logic_vector(to_unsigned(232, 8)),
			1475 => std_logic_vector(to_unsigned(48, 8)),
			1476 => std_logic_vector(to_unsigned(50, 8)),
			1477 => std_logic_vector(to_unsigned(28, 8)),
			1478 => std_logic_vector(to_unsigned(47, 8)),
			1479 => std_logic_vector(to_unsigned(23, 8)),
			1480 => std_logic_vector(to_unsigned(142, 8)),
			1481 => std_logic_vector(to_unsigned(13, 8)),
			1482 => std_logic_vector(to_unsigned(250, 8)),
			1483 => std_logic_vector(to_unsigned(84, 8)),
			1484 => std_logic_vector(to_unsigned(137, 8)),
			1485 => std_logic_vector(to_unsigned(163, 8)),
			1486 => std_logic_vector(to_unsigned(155, 8)),
			1487 => std_logic_vector(to_unsigned(153, 8)),
			1488 => std_logic_vector(to_unsigned(123, 8)),
			1489 => std_logic_vector(to_unsigned(106, 8)),
			1490 => std_logic_vector(to_unsigned(168, 8)),
			1491 => std_logic_vector(to_unsigned(125, 8)),
			1492 => std_logic_vector(to_unsigned(58, 8)),
			1493 => std_logic_vector(to_unsigned(238, 8)),
			1494 => std_logic_vector(to_unsigned(197, 8)),
			1495 => std_logic_vector(to_unsigned(83, 8)),
			1496 => std_logic_vector(to_unsigned(182, 8)),
			1497 => std_logic_vector(to_unsigned(199, 8)),
			1498 => std_logic_vector(to_unsigned(54, 8)),
			1499 => std_logic_vector(to_unsigned(93, 8)),
			1500 => std_logic_vector(to_unsigned(47, 8)),
			1501 => std_logic_vector(to_unsigned(96, 8)),
			1502 => std_logic_vector(to_unsigned(124, 8)),
			1503 => std_logic_vector(to_unsigned(170, 8)),
			1504 => std_logic_vector(to_unsigned(199, 8)),
			1505 => std_logic_vector(to_unsigned(227, 8)),
			1506 => std_logic_vector(to_unsigned(130, 8)),
			1507 => std_logic_vector(to_unsigned(68, 8)),
			1508 => std_logic_vector(to_unsigned(228, 8)),
			1509 => std_logic_vector(to_unsigned(38, 8)),
			1510 => std_logic_vector(to_unsigned(62, 8)),
			1511 => std_logic_vector(to_unsigned(110, 8)),
			1512 => std_logic_vector(to_unsigned(181, 8)),
			1513 => std_logic_vector(to_unsigned(236, 8)),
			1514 => std_logic_vector(to_unsigned(39, 8)),
			1515 => std_logic_vector(to_unsigned(36, 8)),
			1516 => std_logic_vector(to_unsigned(158, 8)),
			1517 => std_logic_vector(to_unsigned(108, 8)),
			1518 => std_logic_vector(to_unsigned(164, 8)),
			1519 => std_logic_vector(to_unsigned(145, 8)),
			1520 => std_logic_vector(to_unsigned(59, 8)),
			1521 => std_logic_vector(to_unsigned(162, 8)),
			1522 => std_logic_vector(to_unsigned(174, 8)),
			1523 => std_logic_vector(to_unsigned(64, 8)),
			1524 => std_logic_vector(to_unsigned(33, 8)),
			1525 => std_logic_vector(to_unsigned(207, 8)),
			1526 => std_logic_vector(to_unsigned(134, 8)),
			1527 => std_logic_vector(to_unsigned(8, 8)),
			1528 => std_logic_vector(to_unsigned(224, 8)),
			1529 => std_logic_vector(to_unsigned(215, 8)),
			1530 => std_logic_vector(to_unsigned(185, 8)),
			1531 => std_logic_vector(to_unsigned(159, 8)),
			1532 => std_logic_vector(to_unsigned(141, 8)),
			1533 => std_logic_vector(to_unsigned(51, 8)),
			1534 => std_logic_vector(to_unsigned(136, 8)),
			1535 => std_logic_vector(to_unsigned(169, 8)),
			1536 => std_logic_vector(to_unsigned(171, 8)),
			1537 => std_logic_vector(to_unsigned(133, 8)),
			1538 => std_logic_vector(to_unsigned(17, 8)),
			1539 => std_logic_vector(to_unsigned(182, 8)),
			1540 => std_logic_vector(to_unsigned(109, 8)),
			1541 => std_logic_vector(to_unsigned(196, 8)),
			1542 => std_logic_vector(to_unsigned(36, 8)),
			1543 => std_logic_vector(to_unsigned(188, 8)),
			1544 => std_logic_vector(to_unsigned(61, 8)),
			1545 => std_logic_vector(to_unsigned(214, 8)),
			1546 => std_logic_vector(to_unsigned(213, 8)),
			1547 => std_logic_vector(to_unsigned(221, 8)),
			1548 => std_logic_vector(to_unsigned(223, 8)),
			1549 => std_logic_vector(to_unsigned(201, 8)),
			1550 => std_logic_vector(to_unsigned(66, 8)),
			1551 => std_logic_vector(to_unsigned(71, 8)),
			1552 => std_logic_vector(to_unsigned(80, 8)),
			1553 => std_logic_vector(to_unsigned(137, 8)),
			1554 => std_logic_vector(to_unsigned(65, 8)),
			1555 => std_logic_vector(to_unsigned(202, 8)),
			1556 => std_logic_vector(to_unsigned(37, 8)),
			1557 => std_logic_vector(to_unsigned(179, 8)),
			1558 => std_logic_vector(to_unsigned(101, 8)),
			1559 => std_logic_vector(to_unsigned(0, 8)),
			1560 => std_logic_vector(to_unsigned(201, 8)),
			1561 => std_logic_vector(to_unsigned(57, 8)),
			1562 => std_logic_vector(to_unsigned(96, 8)),
			1563 => std_logic_vector(to_unsigned(122, 8)),
			1564 => std_logic_vector(to_unsigned(179, 8)),
			1565 => std_logic_vector(to_unsigned(91, 8)),
			1566 => std_logic_vector(to_unsigned(245, 8)),
			1567 => std_logic_vector(to_unsigned(175, 8)),
			1568 => std_logic_vector(to_unsigned(37, 8)),
			1569 => std_logic_vector(to_unsigned(93, 8)),
			1570 => std_logic_vector(to_unsigned(39, 8)),
			1571 => std_logic_vector(to_unsigned(160, 8)),
			1572 => std_logic_vector(to_unsigned(147, 8)),
			1573 => std_logic_vector(to_unsigned(119, 8)),
			1574 => std_logic_vector(to_unsigned(22, 8)),
			1575 => std_logic_vector(to_unsigned(154, 8)),
			1576 => std_logic_vector(to_unsigned(14, 8)),
			1577 => std_logic_vector(to_unsigned(105, 8)),
			1578 => std_logic_vector(to_unsigned(97, 8)),
			1579 => std_logic_vector(to_unsigned(174, 8)),
			1580 => std_logic_vector(to_unsigned(215, 8)),
			1581 => std_logic_vector(to_unsigned(113, 8)),
			1582 => std_logic_vector(to_unsigned(126, 8)),
			1583 => std_logic_vector(to_unsigned(7, 8)),
			1584 => std_logic_vector(to_unsigned(231, 8)),
			1585 => std_logic_vector(to_unsigned(92, 8)),
			1586 => std_logic_vector(to_unsigned(196, 8)),
			1587 => std_logic_vector(to_unsigned(147, 8)),
			1588 => std_logic_vector(to_unsigned(229, 8)),
			1589 => std_logic_vector(to_unsigned(94, 8)),
			1590 => std_logic_vector(to_unsigned(8, 8)),
			1591 => std_logic_vector(to_unsigned(248, 8)),
			1592 => std_logic_vector(to_unsigned(161, 8)),
			1593 => std_logic_vector(to_unsigned(59, 8)),
			1594 => std_logic_vector(to_unsigned(10, 8)),
			1595 => std_logic_vector(to_unsigned(1, 8)),
			1596 => std_logic_vector(to_unsigned(164, 8)),
			1597 => std_logic_vector(to_unsigned(117, 8)),
			1598 => std_logic_vector(to_unsigned(202, 8)),
			1599 => std_logic_vector(to_unsigned(40, 8)),
			1600 => std_logic_vector(to_unsigned(202, 8)),
			1601 => std_logic_vector(to_unsigned(163, 8)),
			1602 => std_logic_vector(to_unsigned(58, 8)),
			1603 => std_logic_vector(to_unsigned(199, 8)),
			1604 => std_logic_vector(to_unsigned(236, 8)),
			1605 => std_logic_vector(to_unsigned(25, 8)),
			1606 => std_logic_vector(to_unsigned(225, 8)),
			1607 => std_logic_vector(to_unsigned(134, 8)),
			1608 => std_logic_vector(to_unsigned(176, 8)),
			1609 => std_logic_vector(to_unsigned(209, 8)),
			1610 => std_logic_vector(to_unsigned(6, 8)),
			1611 => std_logic_vector(to_unsigned(25, 8)),
			1612 => std_logic_vector(to_unsigned(252, 8)),
			1613 => std_logic_vector(to_unsigned(163, 8)),
			1614 => std_logic_vector(to_unsigned(42, 8)),
			1615 => std_logic_vector(to_unsigned(249, 8)),
			1616 => std_logic_vector(to_unsigned(136, 8)),
			1617 => std_logic_vector(to_unsigned(235, 8)),
			1618 => std_logic_vector(to_unsigned(172, 8)),
			1619 => std_logic_vector(to_unsigned(128, 8)),
			1620 => std_logic_vector(to_unsigned(61, 8)),
			1621 => std_logic_vector(to_unsigned(185, 8)),
			1622 => std_logic_vector(to_unsigned(114, 8)),
			1623 => std_logic_vector(to_unsigned(163, 8)),
			1624 => std_logic_vector(to_unsigned(204, 8)),
			1625 => std_logic_vector(to_unsigned(5, 8)),
			1626 => std_logic_vector(to_unsigned(150, 8)),
			1627 => std_logic_vector(to_unsigned(22, 8)),
			1628 => std_logic_vector(to_unsigned(22, 8)),
			1629 => std_logic_vector(to_unsigned(157, 8)),
			1630 => std_logic_vector(to_unsigned(46, 8)),
			1631 => std_logic_vector(to_unsigned(220, 8)),
			1632 => std_logic_vector(to_unsigned(160, 8)),
			1633 => std_logic_vector(to_unsigned(72, 8)),
			1634 => std_logic_vector(to_unsigned(202, 8)),
			1635 => std_logic_vector(to_unsigned(82, 8)),
			1636 => std_logic_vector(to_unsigned(254, 8)),
			1637 => std_logic_vector(to_unsigned(242, 8)),
			1638 => std_logic_vector(to_unsigned(172, 8)),
			1639 => std_logic_vector(to_unsigned(141, 8)),
			1640 => std_logic_vector(to_unsigned(80, 8)),
			1641 => std_logic_vector(to_unsigned(222, 8)),
			1642 => std_logic_vector(to_unsigned(72, 8)),
			1643 => std_logic_vector(to_unsigned(189, 8)),
			1644 => std_logic_vector(to_unsigned(177, 8)),
			1645 => std_logic_vector(to_unsigned(54, 8)),
			1646 => std_logic_vector(to_unsigned(67, 8)),
			1647 => std_logic_vector(to_unsigned(251, 8)),
			1648 => std_logic_vector(to_unsigned(84, 8)),
			1649 => std_logic_vector(to_unsigned(37, 8)),
			1650 => std_logic_vector(to_unsigned(246, 8)),
			1651 => std_logic_vector(to_unsigned(238, 8)),
			1652 => std_logic_vector(to_unsigned(64, 8)),
			1653 => std_logic_vector(to_unsigned(150, 8)),
			1654 => std_logic_vector(to_unsigned(64, 8)),
			1655 => std_logic_vector(to_unsigned(21, 8)),
			1656 => std_logic_vector(to_unsigned(18, 8)),
			1657 => std_logic_vector(to_unsigned(33, 8)),
			others => (others => '0'));             

component project_reti_logiche is
port (
      i_clk         : in  std_logic;
      i_start       : in  std_logic;
      i_rst         : in  std_logic;
      i_data        : in  std_logic_vector(7 downto 0);
      o_address     : out std_logic_vector(15 downto 0);
      o_done        : out std_logic;
      o_en          : out std_logic;
      o_we          : out std_logic;
      o_data        : out std_logic_vector (7 downto 0)
      );
end component project_reti_logiche;


begin
UUT: project_reti_logiche
port map (
          i_clk      	=> tb_clk,
          i_start       => tb_start,
          i_rst      	=> tb_rst,
          i_data    	=> mem_o_data,
          o_address  	=> mem_address,
          o_done      	=> tb_done,
          o_en   	=> enable_wire,
          o_we 		=> mem_we,
          o_data    	=> mem_i_data
          );

p_CLK_GEN : process is
begin
    wait for c_CLOCK_PERIOD/2;
    tb_clk <= not tb_clk;
end process p_CLK_GEN;


MEM : process(tb_clk)
begin
if tb_clk'event and tb_clk = '1' then
    if enable_wire = '1' then
        if i = "00" then
            if mem_we = '1' then
                RAM(conv_integer(mem_address))  <= mem_i_data;
                mem_o_data                      <= mem_i_data after 1 ns;
            else
                mem_o_data <= RAM(conv_integer(mem_address)) after 1 ns;
            end if;
        elsif i ="01" then
            if mem_we = '1' then
                RAM1(conv_integer(mem_address))  <= mem_i_data;
                mem_o_data                      <= mem_i_data after 1 ns;
            else
                mem_o_data <= RAM1(conv_integer(mem_address)) after 1 ns;
            end if;
        elsif i = "10" then 
            if mem_we = '1' then
                RAM2(conv_integer(mem_address))  <= mem_i_data;
                mem_o_data                      <= mem_i_data after 1 ns;
            else
                mem_o_data <= RAM2(conv_integer(mem_address)) after 1 ns;
            end if;
        end if;
    end if;
end if;
end process;


test : process is
begin 
    wait for 100 ns;
    wait for c_CLOCK_PERIOD;
    tb_rst <= '1';
    wait for c_CLOCK_PERIOD;
    wait for 100 ns;
    tb_rst <= '0';
    wait for c_CLOCK_PERIOD;
    wait for 100 ns;
    tb_start <= '1';
    wait for c_CLOCK_PERIOD*75;
	tb_start <= '0';
	tb_rst <= '1';
	wait for c_CLOCK_PERIOD;
	tb_rst <= '0';
	tb_start <= '1';
    wait until tb_done = '1';
    wait for c_CLOCK_PERIOD;
    tb_start <= '0';
    wait until tb_done = '0';
    wait for 100 ns;
    i <= "01";

    
    wait for 100 ns;
    tb_start <= '1';
    wait for c_CLOCK_PERIOD;
    wait until tb_done = '1';
    wait for c_CLOCK_PERIOD;
    tb_start <= '0';
    wait until tb_done = '0';
    wait for 100 ns;
    i <= "10";

    
    wait for 100 ns;
    tb_start <= '1';
    wait for c_CLOCK_PERIOD;
    wait until tb_done = '1';
    wait for c_CLOCK_PERIOD;
    tb_start <= '0';
    wait until tb_done = '0';
    wait for 100 ns;
    
	assert RAM(1724) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(1724))))  severity failure;
	assert RAM(1725) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(1725))))  severity failure;
	assert RAM(1726) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(1726))))  severity failure;
	assert RAM(1727) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(1727))))  severity failure;
	assert RAM(1728) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(1728))))  severity failure;
	assert RAM(1729) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(1729))))  severity failure;
	assert RAM(1730) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(1730))))  severity failure;
	assert RAM(1731) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(1731))))  severity failure;
	assert RAM(1732) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(1732))))  severity failure;
	assert RAM(1733) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(1733))))  severity failure;
	assert RAM(1734) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(1734))))  severity failure;
	assert RAM(1735) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(1735))))  severity failure;
	assert RAM(1736) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(1736))))  severity failure;
	assert RAM(1737) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(1737))))  severity failure;
	assert RAM(1738) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(1738))))  severity failure;
	assert RAM(1739) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(1739))))  severity failure;
	assert RAM(1740) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(1740))))  severity failure;
	assert RAM(1741) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(1741))))  severity failure;
	assert RAM(1742) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(1742))))  severity failure;
	assert RAM(1743) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(1743))))  severity failure;
	assert RAM(1744) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(1744))))  severity failure;
	assert RAM(1745) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(1745))))  severity failure;
	assert RAM(1746) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(1746))))  severity failure;
	assert RAM(1747) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(1747))))  severity failure;
	assert RAM(1748) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(1748))))  severity failure;
	assert RAM(1749) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(1749))))  severity failure;
	assert RAM(1750) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(1750))))  severity failure;
	assert RAM(1751) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(1751))))  severity failure;
	assert RAM(1752) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(1752))))  severity failure;
	assert RAM(1753) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(1753))))  severity failure;
	assert RAM(1754) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(1754))))  severity failure;
	assert RAM(1755) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(1755))))  severity failure;
	assert RAM(1756) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(1756))))  severity failure;
	assert RAM(1757) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(1757))))  severity failure;
	assert RAM(1758) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(1758))))  severity failure;
	assert RAM(1759) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(1759))))  severity failure;
	assert RAM(1760) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(1760))))  severity failure;
	assert RAM(1761) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(1761))))  severity failure;
	assert RAM(1762) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(1762))))  severity failure;
	assert RAM(1763) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(1763))))  severity failure;
	assert RAM(1764) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(1764))))  severity failure;
	assert RAM(1765) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(1765))))  severity failure;
	assert RAM(1766) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(1766))))  severity failure;
	assert RAM(1767) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(1767))))  severity failure;
	assert RAM(1768) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(1768))))  severity failure;
	assert RAM(1769) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(1769))))  severity failure;
	assert RAM(1770) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(1770))))  severity failure;
	assert RAM(1771) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(1771))))  severity failure;
	assert RAM(1772) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(1772))))  severity failure;
	assert RAM(1773) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(1773))))  severity failure;
	assert RAM(1774) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(1774))))  severity failure;
	assert RAM(1775) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(1775))))  severity failure;
	assert RAM(1776) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(1776))))  severity failure;
	assert RAM(1777) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(1777))))  severity failure;
	assert RAM(1778) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(1778))))  severity failure;
	assert RAM(1779) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(1779))))  severity failure;
	assert RAM(1780) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(1780))))  severity failure;
	assert RAM(1781) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(1781))))  severity failure;
	assert RAM(1782) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(1782))))  severity failure;
	assert RAM(1783) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(1783))))  severity failure;
	assert RAM(1784) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(1784))))  severity failure;
	assert RAM(1785) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(1785))))  severity failure;
	assert RAM(1786) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(1786))))  severity failure;
	assert RAM(1787) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(1787))))  severity failure;
	assert RAM(1788) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(1788))))  severity failure;
	assert RAM(1789) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(1789))))  severity failure;
	assert RAM(1790) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(1790))))  severity failure;
	assert RAM(1791) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(1791))))  severity failure;
	assert RAM(1792) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(1792))))  severity failure;
	assert RAM(1793) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(1793))))  severity failure;
	assert RAM(1794) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(1794))))  severity failure;
	assert RAM(1795) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(1795))))  severity failure;
	assert RAM(1796) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(1796))))  severity failure;
	assert RAM(1797) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(1797))))  severity failure;
	assert RAM(1798) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(1798))))  severity failure;
	assert RAM(1799) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(1799))))  severity failure;
	assert RAM(1800) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(1800))))  severity failure;
	assert RAM(1801) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(1801))))  severity failure;
	assert RAM(1802) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(1802))))  severity failure;
	assert RAM(1803) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(1803))))  severity failure;
	assert RAM(1804) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(1804))))  severity failure;
	assert RAM(1805) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(1805))))  severity failure;
	assert RAM(1806) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(1806))))  severity failure;
	assert RAM(1807) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(1807))))  severity failure;
	assert RAM(1808) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(1808))))  severity failure;
	assert RAM(1809) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(1809))))  severity failure;
	assert RAM(1810) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(1810))))  severity failure;
	assert RAM(1811) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(1811))))  severity failure;
	assert RAM(1812) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(1812))))  severity failure;
	assert RAM(1813) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(1813))))  severity failure;
	assert RAM(1814) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(1814))))  severity failure;
	assert RAM(1815) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(1815))))  severity failure;
	assert RAM(1816) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(1816))))  severity failure;
	assert RAM(1817) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(1817))))  severity failure;
	assert RAM(1818) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(1818))))  severity failure;
	assert RAM(1819) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(1819))))  severity failure;
	assert RAM(1820) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(1820))))  severity failure;
	assert RAM(1821) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(1821))))  severity failure;
	assert RAM(1822) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(1822))))  severity failure;
	assert RAM(1823) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(1823))))  severity failure;
	assert RAM(1824) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(1824))))  severity failure;
	assert RAM(1825) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(1825))))  severity failure;
	assert RAM(1826) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(1826))))  severity failure;
	assert RAM(1827) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(1827))))  severity failure;
	assert RAM(1828) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(1828))))  severity failure;
	assert RAM(1829) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(1829))))  severity failure;
	assert RAM(1830) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(1830))))  severity failure;
	assert RAM(1831) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(1831))))  severity failure;
	assert RAM(1832) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(1832))))  severity failure;
	assert RAM(1833) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(1833))))  severity failure;
	assert RAM(1834) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(1834))))  severity failure;
	assert RAM(1835) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(1835))))  severity failure;
	assert RAM(1836) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(1836))))  severity failure;
	assert RAM(1837) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(1837))))  severity failure;
	assert RAM(1838) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(1838))))  severity failure;
	assert RAM(1839) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(1839))))  severity failure;
	assert RAM(1840) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(1840))))  severity failure;
	assert RAM(1841) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(1841))))  severity failure;
	assert RAM(1842) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(1842))))  severity failure;
	assert RAM(1843) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(1843))))  severity failure;
	assert RAM(1844) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(1844))))  severity failure;
	assert RAM(1845) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(1845))))  severity failure;
	assert RAM(1846) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(1846))))  severity failure;
	assert RAM(1847) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(1847))))  severity failure;
	assert RAM(1848) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(1848))))  severity failure;
	assert RAM(1849) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(1849))))  severity failure;
	assert RAM(1850) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(1850))))  severity failure;
	assert RAM(1851) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(1851))))  severity failure;
	assert RAM(1852) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(1852))))  severity failure;
	assert RAM(1853) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(1853))))  severity failure;
	assert RAM(1854) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(1854))))  severity failure;
	assert RAM(1855) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(1855))))  severity failure;
	assert RAM(1856) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(1856))))  severity failure;
	assert RAM(1857) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(1857))))  severity failure;
	assert RAM(1858) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(1858))))  severity failure;
	assert RAM(1859) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(1859))))  severity failure;
	assert RAM(1860) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(1860))))  severity failure;
	assert RAM(1861) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(1861))))  severity failure;
	assert RAM(1862) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(1862))))  severity failure;
	assert RAM(1863) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(1863))))  severity failure;
	assert RAM(1864) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(1864))))  severity failure;
	assert RAM(1865) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(1865))))  severity failure;
	assert RAM(1866) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(1866))))  severity failure;
	assert RAM(1867) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(1867))))  severity failure;
	assert RAM(1868) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(1868))))  severity failure;
	assert RAM(1869) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(1869))))  severity failure;
	assert RAM(1870) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(1870))))  severity failure;
	assert RAM(1871) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(1871))))  severity failure;
	assert RAM(1872) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(1872))))  severity failure;
	assert RAM(1873) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(1873))))  severity failure;
	assert RAM(1874) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(1874))))  severity failure;
	assert RAM(1875) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(1875))))  severity failure;
	assert RAM(1876) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(1876))))  severity failure;
	assert RAM(1877) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(1877))))  severity failure;
	assert RAM(1878) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(1878))))  severity failure;
	assert RAM(1879) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(1879))))  severity failure;
	assert RAM(1880) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(1880))))  severity failure;
	assert RAM(1881) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(1881))))  severity failure;
	assert RAM(1882) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(1882))))  severity failure;
	assert RAM(1883) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(1883))))  severity failure;
	assert RAM(1884) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(1884))))  severity failure;
	assert RAM(1885) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(1885))))  severity failure;
	assert RAM(1886) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(1886))))  severity failure;
	assert RAM(1887) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(1887))))  severity failure;
	assert RAM(1888) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(1888))))  severity failure;
	assert RAM(1889) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(1889))))  severity failure;
	assert RAM(1890) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(1890))))  severity failure;
	assert RAM(1891) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(1891))))  severity failure;
	assert RAM(1892) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(1892))))  severity failure;
	assert RAM(1893) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(1893))))  severity failure;
	assert RAM(1894) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(1894))))  severity failure;
	assert RAM(1895) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(1895))))  severity failure;
	assert RAM(1896) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(1896))))  severity failure;
	assert RAM(1897) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(1897))))  severity failure;
	assert RAM(1898) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(1898))))  severity failure;
	assert RAM(1899) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(1899))))  severity failure;
	assert RAM(1900) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(1900))))  severity failure;
	assert RAM(1901) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(1901))))  severity failure;
	assert RAM(1902) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(1902))))  severity failure;
	assert RAM(1903) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(1903))))  severity failure;
	assert RAM(1904) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(1904))))  severity failure;
	assert RAM(1905) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(1905))))  severity failure;
	assert RAM(1906) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(1906))))  severity failure;
	assert RAM(1907) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(1907))))  severity failure;
	assert RAM(1908) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(1908))))  severity failure;
	assert RAM(1909) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(1909))))  severity failure;
	assert RAM(1910) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(1910))))  severity failure;
	assert RAM(1911) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(1911))))  severity failure;
	assert RAM(1912) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(1912))))  severity failure;
	assert RAM(1913) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(1913))))  severity failure;
	assert RAM(1914) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(1914))))  severity failure;
	assert RAM(1915) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(1915))))  severity failure;
	assert RAM(1916) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(1916))))  severity failure;
	assert RAM(1917) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(1917))))  severity failure;
	assert RAM(1918) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(1918))))  severity failure;
	assert RAM(1919) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(1919))))  severity failure;
	assert RAM(1920) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(1920))))  severity failure;
	assert RAM(1921) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(1921))))  severity failure;
	assert RAM(1922) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(1922))))  severity failure;
	assert RAM(1923) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(1923))))  severity failure;
	assert RAM(1924) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(1924))))  severity failure;
	assert RAM(1925) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(1925))))  severity failure;
	assert RAM(1926) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(1926))))  severity failure;
	assert RAM(1927) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(1927))))  severity failure;
	assert RAM(1928) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(1928))))  severity failure;
	assert RAM(1929) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(1929))))  severity failure;
	assert RAM(1930) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(1930))))  severity failure;
	assert RAM(1931) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(1931))))  severity failure;
	assert RAM(1932) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(1932))))  severity failure;
	assert RAM(1933) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(1933))))  severity failure;
	assert RAM(1934) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(1934))))  severity failure;
	assert RAM(1935) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(1935))))  severity failure;
	assert RAM(1936) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(1936))))  severity failure;
	assert RAM(1937) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(1937))))  severity failure;
	assert RAM(1938) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(1938))))  severity failure;
	assert RAM(1939) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(1939))))  severity failure;
	assert RAM(1940) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(1940))))  severity failure;
	assert RAM(1941) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(1941))))  severity failure;
	assert RAM(1942) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(1942))))  severity failure;
	assert RAM(1943) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(1943))))  severity failure;
	assert RAM(1944) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(1944))))  severity failure;
	assert RAM(1945) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(1945))))  severity failure;
	assert RAM(1946) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(1946))))  severity failure;
	assert RAM(1947) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(1947))))  severity failure;
	assert RAM(1948) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(1948))))  severity failure;
	assert RAM(1949) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(1949))))  severity failure;
	assert RAM(1950) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(1950))))  severity failure;
	assert RAM(1951) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(1951))))  severity failure;
	assert RAM(1952) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(1952))))  severity failure;
	assert RAM(1953) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(1953))))  severity failure;
	assert RAM(1954) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(1954))))  severity failure;
	assert RAM(1955) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(1955))))  severity failure;
	assert RAM(1956) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(1956))))  severity failure;
	assert RAM(1957) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(1957))))  severity failure;
	assert RAM(1958) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(1958))))  severity failure;
	assert RAM(1959) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(1959))))  severity failure;
	assert RAM(1960) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(1960))))  severity failure;
	assert RAM(1961) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(1961))))  severity failure;
	assert RAM(1962) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(1962))))  severity failure;
	assert RAM(1963) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(1963))))  severity failure;
	assert RAM(1964) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(1964))))  severity failure;
	assert RAM(1965) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(1965))))  severity failure;
	assert RAM(1966) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(1966))))  severity failure;
	assert RAM(1967) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(1967))))  severity failure;
	assert RAM(1968) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(1968))))  severity failure;
	assert RAM(1969) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(1969))))  severity failure;
	assert RAM(1970) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(1970))))  severity failure;
	assert RAM(1971) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(1971))))  severity failure;
	assert RAM(1972) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(1972))))  severity failure;
	assert RAM(1973) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(1973))))  severity failure;
	assert RAM(1974) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(1974))))  severity failure;
	assert RAM(1975) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(1975))))  severity failure;
	assert RAM(1976) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(1976))))  severity failure;
	assert RAM(1977) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(1977))))  severity failure;
	assert RAM(1978) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(1978))))  severity failure;
	assert RAM(1979) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(1979))))  severity failure;
	assert RAM(1980) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(1980))))  severity failure;
	assert RAM(1981) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(1981))))  severity failure;
	assert RAM(1982) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(1982))))  severity failure;
	assert RAM(1983) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(1983))))  severity failure;
	assert RAM(1984) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(1984))))  severity failure;
	assert RAM(1985) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(1985))))  severity failure;
	assert RAM(1986) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(1986))))  severity failure;
	assert RAM(1987) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(1987))))  severity failure;
	assert RAM(1988) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(1988))))  severity failure;
	assert RAM(1989) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(1989))))  severity failure;
	assert RAM(1990) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(1990))))  severity failure;
	assert RAM(1991) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(1991))))  severity failure;
	assert RAM(1992) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(1992))))  severity failure;
	assert RAM(1993) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(1993))))  severity failure;
	assert RAM(1994) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(1994))))  severity failure;
	assert RAM(1995) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(1995))))  severity failure;
	assert RAM(1996) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(1996))))  severity failure;
	assert RAM(1997) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(1997))))  severity failure;
	assert RAM(1998) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(1998))))  severity failure;
	assert RAM(1999) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(1999))))  severity failure;
	assert RAM(2000) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(2000))))  severity failure;
	assert RAM(2001) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(2001))))  severity failure;
	assert RAM(2002) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(2002))))  severity failure;
	assert RAM(2003) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(2003))))  severity failure;
	assert RAM(2004) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(2004))))  severity failure;
	assert RAM(2005) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(2005))))  severity failure;
	assert RAM(2006) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(2006))))  severity failure;
	assert RAM(2007) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(2007))))  severity failure;
	assert RAM(2008) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(2008))))  severity failure;
	assert RAM(2009) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(2009))))  severity failure;
	assert RAM(2010) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(2010))))  severity failure;
	assert RAM(2011) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(2011))))  severity failure;
	assert RAM(2012) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(2012))))  severity failure;
	assert RAM(2013) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(2013))))  severity failure;
	assert RAM(2014) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(2014))))  severity failure;
	assert RAM(2015) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(2015))))  severity failure;
	assert RAM(2016) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(2016))))  severity failure;
	assert RAM(2017) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(2017))))  severity failure;
	assert RAM(2018) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(2018))))  severity failure;
	assert RAM(2019) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(2019))))  severity failure;
	assert RAM(2020) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(2020))))  severity failure;
	assert RAM(2021) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(2021))))  severity failure;
	assert RAM(2022) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(2022))))  severity failure;
	assert RAM(2023) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(2023))))  severity failure;
	assert RAM(2024) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(2024))))  severity failure;
	assert RAM(2025) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(2025))))  severity failure;
	assert RAM(2026) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(2026))))  severity failure;
	assert RAM(2027) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(2027))))  severity failure;
	assert RAM(2028) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(2028))))  severity failure;
	assert RAM(2029) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(2029))))  severity failure;
	assert RAM(2030) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(2030))))  severity failure;
	assert RAM(2031) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(2031))))  severity failure;
	assert RAM(2032) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(2032))))  severity failure;
	assert RAM(2033) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(2033))))  severity failure;
	assert RAM(2034) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(2034))))  severity failure;
	assert RAM(2035) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(2035))))  severity failure;
	assert RAM(2036) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(2036))))  severity failure;
	assert RAM(2037) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(2037))))  severity failure;
	assert RAM(2038) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(2038))))  severity failure;
	assert RAM(2039) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(2039))))  severity failure;
	assert RAM(2040) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(2040))))  severity failure;
	assert RAM(2041) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(2041))))  severity failure;
	assert RAM(2042) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(2042))))  severity failure;
	assert RAM(2043) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(2043))))  severity failure;
	assert RAM(2044) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(2044))))  severity failure;
	assert RAM(2045) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(2045))))  severity failure;
	assert RAM(2046) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(2046))))  severity failure;
	assert RAM(2047) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(2047))))  severity failure;
	assert RAM(2048) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(2048))))  severity failure;
	assert RAM(2049) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(2049))))  severity failure;
	assert RAM(2050) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(2050))))  severity failure;
	assert RAM(2051) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(2051))))  severity failure;
	assert RAM(2052) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(2052))))  severity failure;
	assert RAM(2053) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(2053))))  severity failure;
	assert RAM(2054) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(2054))))  severity failure;
	assert RAM(2055) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(2055))))  severity failure;
	assert RAM(2056) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(2056))))  severity failure;
	assert RAM(2057) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(2057))))  severity failure;
	assert RAM(2058) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(2058))))  severity failure;
	assert RAM(2059) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(2059))))  severity failure;
	assert RAM(2060) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(2060))))  severity failure;
	assert RAM(2061) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(2061))))  severity failure;
	assert RAM(2062) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(2062))))  severity failure;
	assert RAM(2063) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(2063))))  severity failure;
	assert RAM(2064) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(2064))))  severity failure;
	assert RAM(2065) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(2065))))  severity failure;
	assert RAM(2066) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(2066))))  severity failure;
	assert RAM(2067) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(2067))))  severity failure;
	assert RAM(2068) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(2068))))  severity failure;
	assert RAM(2069) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(2069))))  severity failure;
	assert RAM(2070) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(2070))))  severity failure;
	assert RAM(2071) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(2071))))  severity failure;
	assert RAM(2072) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(2072))))  severity failure;
	assert RAM(2073) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(2073))))  severity failure;
	assert RAM(2074) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(2074))))  severity failure;
	assert RAM(2075) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(2075))))  severity failure;
	assert RAM(2076) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(2076))))  severity failure;
	assert RAM(2077) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(2077))))  severity failure;
	assert RAM(2078) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(2078))))  severity failure;
	assert RAM(2079) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(2079))))  severity failure;
	assert RAM(2080) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(2080))))  severity failure;
	assert RAM(2081) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(2081))))  severity failure;
	assert RAM(2082) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(2082))))  severity failure;
	assert RAM(2083) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(2083))))  severity failure;
	assert RAM(2084) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(2084))))  severity failure;
	assert RAM(2085) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(2085))))  severity failure;
	assert RAM(2086) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(2086))))  severity failure;
	assert RAM(2087) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(2087))))  severity failure;
	assert RAM(2088) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(2088))))  severity failure;
	assert RAM(2089) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(2089))))  severity failure;
	assert RAM(2090) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(2090))))  severity failure;
	assert RAM(2091) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(2091))))  severity failure;
	assert RAM(2092) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(2092))))  severity failure;
	assert RAM(2093) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(2093))))  severity failure;
	assert RAM(2094) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(2094))))  severity failure;
	assert RAM(2095) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(2095))))  severity failure;
	assert RAM(2096) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(2096))))  severity failure;
	assert RAM(2097) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(2097))))  severity failure;
	assert RAM(2098) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(2098))))  severity failure;
	assert RAM(2099) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(2099))))  severity failure;
	assert RAM(2100) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(2100))))  severity failure;
	assert RAM(2101) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(2101))))  severity failure;
	assert RAM(2102) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(2102))))  severity failure;
	assert RAM(2103) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(2103))))  severity failure;
	assert RAM(2104) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(2104))))  severity failure;
	assert RAM(2105) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(2105))))  severity failure;
	assert RAM(2106) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(2106))))  severity failure;
	assert RAM(2107) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(2107))))  severity failure;
	assert RAM(2108) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(2108))))  severity failure;
	assert RAM(2109) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(2109))))  severity failure;
	assert RAM(2110) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(2110))))  severity failure;
	assert RAM(2111) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(2111))))  severity failure;
	assert RAM(2112) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(2112))))  severity failure;
	assert RAM(2113) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(2113))))  severity failure;
	assert RAM(2114) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(2114))))  severity failure;
	assert RAM(2115) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(2115))))  severity failure;
	assert RAM(2116) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(2116))))  severity failure;
	assert RAM(2117) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(2117))))  severity failure;
	assert RAM(2118) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(2118))))  severity failure;
	assert RAM(2119) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(2119))))  severity failure;
	assert RAM(2120) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(2120))))  severity failure;
	assert RAM(2121) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(2121))))  severity failure;
	assert RAM(2122) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(2122))))  severity failure;
	assert RAM(2123) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(2123))))  severity failure;
	assert RAM(2124) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(2124))))  severity failure;
	assert RAM(2125) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(2125))))  severity failure;
	assert RAM(2126) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(2126))))  severity failure;
	assert RAM(2127) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(2127))))  severity failure;
	assert RAM(2128) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(2128))))  severity failure;
	assert RAM(2129) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(2129))))  severity failure;
	assert RAM(2130) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(2130))))  severity failure;
	assert RAM(2131) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(2131))))  severity failure;
	assert RAM(2132) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(2132))))  severity failure;
	assert RAM(2133) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(2133))))  severity failure;
	assert RAM(2134) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(2134))))  severity failure;
	assert RAM(2135) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(2135))))  severity failure;
	assert RAM(2136) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(2136))))  severity failure;
	assert RAM(2137) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(2137))))  severity failure;
	assert RAM(2138) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(2138))))  severity failure;
	assert RAM(2139) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(2139))))  severity failure;
	assert RAM(2140) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(2140))))  severity failure;
	assert RAM(2141) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(2141))))  severity failure;
	assert RAM(2142) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(2142))))  severity failure;
	assert RAM(2143) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(2143))))  severity failure;
	assert RAM(2144) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(2144))))  severity failure;
	assert RAM(2145) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(2145))))  severity failure;
	assert RAM(2146) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(2146))))  severity failure;
	assert RAM(2147) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(2147))))  severity failure;
	assert RAM(2148) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(2148))))  severity failure;
	assert RAM(2149) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(2149))))  severity failure;
	assert RAM(2150) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(2150))))  severity failure;
	assert RAM(2151) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(2151))))  severity failure;
	assert RAM(2152) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(2152))))  severity failure;
	assert RAM(2153) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(2153))))  severity failure;
	assert RAM(2154) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(2154))))  severity failure;
	assert RAM(2155) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(2155))))  severity failure;
	assert RAM(2156) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(2156))))  severity failure;
	assert RAM(2157) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(2157))))  severity failure;
	assert RAM(2158) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(2158))))  severity failure;
	assert RAM(2159) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(2159))))  severity failure;
	assert RAM(2160) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(2160))))  severity failure;
	assert RAM(2161) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(2161))))  severity failure;
	assert RAM(2162) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(2162))))  severity failure;
	assert RAM(2163) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(2163))))  severity failure;
	assert RAM(2164) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(2164))))  severity failure;
	assert RAM(2165) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(2165))))  severity failure;
	assert RAM(2166) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(2166))))  severity failure;
	assert RAM(2167) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(2167))))  severity failure;
	assert RAM(2168) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(2168))))  severity failure;
	assert RAM(2169) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(2169))))  severity failure;
	assert RAM(2170) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(2170))))  severity failure;
	assert RAM(2171) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(2171))))  severity failure;
	assert RAM(2172) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(2172))))  severity failure;
	assert RAM(2173) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(2173))))  severity failure;
	assert RAM(2174) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(2174))))  severity failure;
	assert RAM(2175) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(2175))))  severity failure;
	assert RAM(2176) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(2176))))  severity failure;
	assert RAM(2177) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(2177))))  severity failure;
	assert RAM(2178) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(2178))))  severity failure;
	assert RAM(2179) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(2179))))  severity failure;
	assert RAM(2180) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(2180))))  severity failure;
	assert RAM(2181) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(2181))))  severity failure;
	assert RAM(2182) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(2182))))  severity failure;
	assert RAM(2183) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(2183))))  severity failure;
	assert RAM(2184) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(2184))))  severity failure;
	assert RAM(2185) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(2185))))  severity failure;
	assert RAM(2186) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(2186))))  severity failure;
	assert RAM(2187) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(2187))))  severity failure;
	assert RAM(2188) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(2188))))  severity failure;
	assert RAM(2189) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(2189))))  severity failure;
	assert RAM(2190) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(2190))))  severity failure;
	assert RAM(2191) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(2191))))  severity failure;
	assert RAM(2192) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(2192))))  severity failure;
	assert RAM(2193) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(2193))))  severity failure;
	assert RAM(2194) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(2194))))  severity failure;
	assert RAM(2195) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(2195))))  severity failure;
	assert RAM(2196) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(2196))))  severity failure;
	assert RAM(2197) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(2197))))  severity failure;
	assert RAM(2198) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(2198))))  severity failure;
	assert RAM(2199) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(2199))))  severity failure;
	assert RAM(2200) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(2200))))  severity failure;
	assert RAM(2201) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(2201))))  severity failure;
	assert RAM(2202) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(2202))))  severity failure;
	assert RAM(2203) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(2203))))  severity failure;
	assert RAM(2204) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(2204))))  severity failure;
	assert RAM(2205) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(2205))))  severity failure;
	assert RAM(2206) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(2206))))  severity failure;
	assert RAM(2207) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(2207))))  severity failure;
	assert RAM(2208) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(2208))))  severity failure;
	assert RAM(2209) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(2209))))  severity failure;
	assert RAM(2210) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(2210))))  severity failure;
	assert RAM(2211) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(2211))))  severity failure;
	assert RAM(2212) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(2212))))  severity failure;
	assert RAM(2213) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(2213))))  severity failure;
	assert RAM(2214) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(2214))))  severity failure;
	assert RAM(2215) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(2215))))  severity failure;
	assert RAM(2216) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(2216))))  severity failure;
	assert RAM(2217) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(2217))))  severity failure;
	assert RAM(2218) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(2218))))  severity failure;
	assert RAM(2219) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(2219))))  severity failure;
	assert RAM(2220) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(2220))))  severity failure;
	assert RAM(2221) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(2221))))  severity failure;
	assert RAM(2222) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(2222))))  severity failure;
	assert RAM(2223) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(2223))))  severity failure;
	assert RAM(2224) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(2224))))  severity failure;
	assert RAM(2225) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(2225))))  severity failure;
	assert RAM(2226) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(2226))))  severity failure;
	assert RAM(2227) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(2227))))  severity failure;
	assert RAM(2228) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(2228))))  severity failure;
	assert RAM(2229) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(2229))))  severity failure;
	assert RAM(2230) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(2230))))  severity failure;
	assert RAM(2231) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(2231))))  severity failure;
	assert RAM(2232) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(2232))))  severity failure;
	assert RAM(2233) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(2233))))  severity failure;
	assert RAM(2234) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(2234))))  severity failure;
	assert RAM(2235) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(2235))))  severity failure;
	assert RAM(2236) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(2236))))  severity failure;
	assert RAM(2237) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(2237))))  severity failure;
	assert RAM(2238) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(2238))))  severity failure;
	assert RAM(2239) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(2239))))  severity failure;
	assert RAM(2240) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(2240))))  severity failure;
	assert RAM(2241) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(2241))))  severity failure;
	assert RAM(2242) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(2242))))  severity failure;
	assert RAM(2243) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(2243))))  severity failure;
	assert RAM(2244) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(2244))))  severity failure;
	assert RAM(2245) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(2245))))  severity failure;
	assert RAM(2246) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(2246))))  severity failure;
	assert RAM(2247) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(2247))))  severity failure;
	assert RAM(2248) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(2248))))  severity failure;
	assert RAM(2249) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(2249))))  severity failure;
	assert RAM(2250) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(2250))))  severity failure;
	assert RAM(2251) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(2251))))  severity failure;
	assert RAM(2252) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(2252))))  severity failure;
	assert RAM(2253) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(2253))))  severity failure;
	assert RAM(2254) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(2254))))  severity failure;
	assert RAM(2255) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(2255))))  severity failure;
	assert RAM(2256) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(2256))))  severity failure;
	assert RAM(2257) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(2257))))  severity failure;
	assert RAM(2258) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(2258))))  severity failure;
	assert RAM(2259) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(2259))))  severity failure;
	assert RAM(2260) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(2260))))  severity failure;
	assert RAM(2261) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(2261))))  severity failure;
	assert RAM(2262) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(2262))))  severity failure;
	assert RAM(2263) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(2263))))  severity failure;
	assert RAM(2264) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(2264))))  severity failure;
	assert RAM(2265) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(2265))))  severity failure;
	assert RAM(2266) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(2266))))  severity failure;
	assert RAM(2267) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(2267))))  severity failure;
	assert RAM(2268) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(2268))))  severity failure;
	assert RAM(2269) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(2269))))  severity failure;
	assert RAM(2270) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(2270))))  severity failure;
	assert RAM(2271) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(2271))))  severity failure;
	assert RAM(2272) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(2272))))  severity failure;
	assert RAM(2273) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(2273))))  severity failure;
	assert RAM(2274) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(2274))))  severity failure;
	assert RAM(2275) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(2275))))  severity failure;
	assert RAM(2276) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(2276))))  severity failure;
	assert RAM(2277) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(2277))))  severity failure;
	assert RAM(2278) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(2278))))  severity failure;
	assert RAM(2279) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(2279))))  severity failure;
	assert RAM(2280) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(2280))))  severity failure;
	assert RAM(2281) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(2281))))  severity failure;
	assert RAM(2282) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(2282))))  severity failure;
	assert RAM(2283) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(2283))))  severity failure;
	assert RAM(2284) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(2284))))  severity failure;
	assert RAM(2285) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(2285))))  severity failure;
	assert RAM(2286) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(2286))))  severity failure;
	assert RAM(2287) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(2287))))  severity failure;
	assert RAM(2288) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(2288))))  severity failure;
	assert RAM(2289) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(2289))))  severity failure;
	assert RAM(2290) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(2290))))  severity failure;
	assert RAM(2291) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(2291))))  severity failure;
	assert RAM(2292) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(2292))))  severity failure;
	assert RAM(2293) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(2293))))  severity failure;
	assert RAM(2294) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(2294))))  severity failure;
	assert RAM(2295) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(2295))))  severity failure;
	assert RAM(2296) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(2296))))  severity failure;
	assert RAM(2297) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(2297))))  severity failure;
	assert RAM(2298) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(2298))))  severity failure;
	assert RAM(2299) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(2299))))  severity failure;
	assert RAM(2300) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(2300))))  severity failure;
	assert RAM(2301) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(2301))))  severity failure;
	assert RAM(2302) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(2302))))  severity failure;
	assert RAM(2303) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(2303))))  severity failure;
	assert RAM(2304) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(2304))))  severity failure;
	assert RAM(2305) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(2305))))  severity failure;
	assert RAM(2306) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(2306))))  severity failure;
	assert RAM(2307) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(2307))))  severity failure;
	assert RAM(2308) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(2308))))  severity failure;
	assert RAM(2309) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(2309))))  severity failure;
	assert RAM(2310) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(2310))))  severity failure;
	assert RAM(2311) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(2311))))  severity failure;
	assert RAM(2312) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(2312))))  severity failure;
	assert RAM(2313) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(2313))))  severity failure;
	assert RAM(2314) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(2314))))  severity failure;
	assert RAM(2315) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(2315))))  severity failure;
	assert RAM(2316) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(2316))))  severity failure;
	assert RAM(2317) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(2317))))  severity failure;
	assert RAM(2318) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(2318))))  severity failure;
	assert RAM(2319) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(2319))))  severity failure;
	assert RAM(2320) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(2320))))  severity failure;
	assert RAM(2321) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(2321))))  severity failure;
	assert RAM(2322) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(2322))))  severity failure;
	assert RAM(2323) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(2323))))  severity failure;
	assert RAM(2324) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(2324))))  severity failure;
	assert RAM(2325) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(2325))))  severity failure;
	assert RAM(2326) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(2326))))  severity failure;
	assert RAM(2327) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(2327))))  severity failure;
	assert RAM(2328) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(2328))))  severity failure;
	assert RAM(2329) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(2329))))  severity failure;
	assert RAM(2330) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(2330))))  severity failure;
	assert RAM(2331) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(2331))))  severity failure;
	assert RAM(2332) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(2332))))  severity failure;
	assert RAM(2333) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(2333))))  severity failure;
	assert RAM(2334) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(2334))))  severity failure;
	assert RAM(2335) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(2335))))  severity failure;
	assert RAM(2336) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(2336))))  severity failure;
	assert RAM(2337) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(2337))))  severity failure;
	assert RAM(2338) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(2338))))  severity failure;
	assert RAM(2339) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(2339))))  severity failure;
	assert RAM(2340) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(2340))))  severity failure;
	assert RAM(2341) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(2341))))  severity failure;
	assert RAM(2342) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(2342))))  severity failure;
	assert RAM(2343) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(2343))))  severity failure;
	assert RAM(2344) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(2344))))  severity failure;
	assert RAM(2345) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(2345))))  severity failure;
	assert RAM(2346) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(2346))))  severity failure;
	assert RAM(2347) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(2347))))  severity failure;
	assert RAM(2348) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(2348))))  severity failure;
	assert RAM(2349) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(2349))))  severity failure;
	assert RAM(2350) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(2350))))  severity failure;
	assert RAM(2351) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(2351))))  severity failure;
	assert RAM(2352) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(2352))))  severity failure;
	assert RAM(2353) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(2353))))  severity failure;
	assert RAM(2354) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(2354))))  severity failure;
	assert RAM(2355) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(2355))))  severity failure;
	assert RAM(2356) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(2356))))  severity failure;
	assert RAM(2357) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(2357))))  severity failure;
	assert RAM(2358) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(2358))))  severity failure;
	assert RAM(2359) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(2359))))  severity failure;
	assert RAM(2360) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(2360))))  severity failure;
	assert RAM(2361) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(2361))))  severity failure;
	assert RAM(2362) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(2362))))  severity failure;
	assert RAM(2363) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(2363))))  severity failure;
	assert RAM(2364) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(2364))))  severity failure;
	assert RAM(2365) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(2365))))  severity failure;
	assert RAM(2366) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(2366))))  severity failure;
	assert RAM(2367) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(2367))))  severity failure;
	assert RAM(2368) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(2368))))  severity failure;
	assert RAM(2369) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(2369))))  severity failure;
	assert RAM(2370) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(2370))))  severity failure;
	assert RAM(2371) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(2371))))  severity failure;
	assert RAM(2372) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(2372))))  severity failure;
	assert RAM(2373) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(2373))))  severity failure;
	assert RAM(2374) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(2374))))  severity failure;
	assert RAM(2375) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(2375))))  severity failure;
	assert RAM(2376) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(2376))))  severity failure;
	assert RAM(2377) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(2377))))  severity failure;
	assert RAM(2378) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(2378))))  severity failure;
	assert RAM(2379) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(2379))))  severity failure;
	assert RAM(2380) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(2380))))  severity failure;
	assert RAM(2381) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(2381))))  severity failure;
	assert RAM(2382) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(2382))))  severity failure;
	assert RAM(2383) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(2383))))  severity failure;
	assert RAM(2384) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(2384))))  severity failure;
	assert RAM(2385) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(2385))))  severity failure;
	assert RAM(2386) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(2386))))  severity failure;
	assert RAM(2387) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(2387))))  severity failure;
	assert RAM(2388) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(2388))))  severity failure;
	assert RAM(2389) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(2389))))  severity failure;
	assert RAM(2390) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(2390))))  severity failure;
	assert RAM(2391) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(2391))))  severity failure;
	assert RAM(2392) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(2392))))  severity failure;
	assert RAM(2393) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(2393))))  severity failure;
	assert RAM(2394) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(2394))))  severity failure;
	assert RAM(2395) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(2395))))  severity failure;
	assert RAM(2396) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(2396))))  severity failure;
	assert RAM(2397) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(2397))))  severity failure;
	assert RAM(2398) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(2398))))  severity failure;
	assert RAM(2399) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(2399))))  severity failure;
	assert RAM(2400) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(2400))))  severity failure;
	assert RAM(2401) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(2401))))  severity failure;
	assert RAM(2402) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(2402))))  severity failure;
	assert RAM(2403) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(2403))))  severity failure;
	assert RAM(2404) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(2404))))  severity failure;
	assert RAM(2405) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(2405))))  severity failure;
	assert RAM(2406) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(2406))))  severity failure;
	assert RAM(2407) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(2407))))  severity failure;
	assert RAM(2408) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(2408))))  severity failure;
	assert RAM(2409) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(2409))))  severity failure;
	assert RAM(2410) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(2410))))  severity failure;
	assert RAM(2411) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(2411))))  severity failure;
	assert RAM(2412) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(2412))))  severity failure;
	assert RAM(2413) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(2413))))  severity failure;
	assert RAM(2414) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(2414))))  severity failure;
	assert RAM(2415) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(2415))))  severity failure;
	assert RAM(2416) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(2416))))  severity failure;
	assert RAM(2417) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(2417))))  severity failure;
	assert RAM(2418) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(2418))))  severity failure;
	assert RAM(2419) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(2419))))  severity failure;
	assert RAM(2420) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(2420))))  severity failure;
	assert RAM(2421) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(2421))))  severity failure;
	assert RAM(2422) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(2422))))  severity failure;
	assert RAM(2423) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(2423))))  severity failure;
	assert RAM(2424) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(2424))))  severity failure;
	assert RAM(2425) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(2425))))  severity failure;
	assert RAM(2426) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(2426))))  severity failure;
	assert RAM(2427) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(2427))))  severity failure;
	assert RAM(2428) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(2428))))  severity failure;
	assert RAM(2429) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(2429))))  severity failure;
	assert RAM(2430) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(2430))))  severity failure;
	assert RAM(2431) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(2431))))  severity failure;
	assert RAM(2432) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(2432))))  severity failure;
	assert RAM(2433) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(2433))))  severity failure;
	assert RAM(2434) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(2434))))  severity failure;
	assert RAM(2435) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(2435))))  severity failure;
	assert RAM(2436) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(2436))))  severity failure;
	assert RAM(2437) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(2437))))  severity failure;
	assert RAM(2438) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(2438))))  severity failure;
	assert RAM(2439) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(2439))))  severity failure;
	assert RAM(2440) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(2440))))  severity failure;
	assert RAM(2441) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(2441))))  severity failure;
	assert RAM(2442) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(2442))))  severity failure;
	assert RAM(2443) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(2443))))  severity failure;
	assert RAM(2444) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(2444))))  severity failure;
	assert RAM(2445) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(2445))))  severity failure;
	assert RAM(2446) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(2446))))  severity failure;
	assert RAM(2447) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(2447))))  severity failure;
	assert RAM(2448) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(2448))))  severity failure;
	assert RAM(2449) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(2449))))  severity failure;
	assert RAM(2450) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(2450))))  severity failure;
	assert RAM(2451) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(2451))))  severity failure;
	assert RAM(2452) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(2452))))  severity failure;
	assert RAM(2453) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(2453))))  severity failure;
	assert RAM(2454) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(2454))))  severity failure;
	assert RAM(2455) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(2455))))  severity failure;
	assert RAM(2456) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(2456))))  severity failure;
	assert RAM(2457) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(2457))))  severity failure;
	assert RAM(2458) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(2458))))  severity failure;
	assert RAM(2459) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(2459))))  severity failure;
	assert RAM(2460) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(2460))))  severity failure;
	assert RAM(2461) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(2461))))  severity failure;
	assert RAM(2462) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(2462))))  severity failure;
	assert RAM(2463) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(2463))))  severity failure;
	assert RAM(2464) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(2464))))  severity failure;
	assert RAM(2465) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(2465))))  severity failure;
	assert RAM(2466) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(2466))))  severity failure;
	assert RAM(2467) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(2467))))  severity failure;
	assert RAM(2468) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(2468))))  severity failure;
	assert RAM(2469) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(2469))))  severity failure;
	assert RAM(2470) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(2470))))  severity failure;
	assert RAM(2471) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(2471))))  severity failure;
	assert RAM(2472) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(2472))))  severity failure;
	assert RAM(2473) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(2473))))  severity failure;
	assert RAM(2474) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(2474))))  severity failure;
	assert RAM(2475) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(2475))))  severity failure;
	assert RAM(2476) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(2476))))  severity failure;
	assert RAM(2477) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(2477))))  severity failure;
	assert RAM(2478) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(2478))))  severity failure;
	assert RAM(2479) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(2479))))  severity failure;
	assert RAM(2480) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(2480))))  severity failure;
	assert RAM(2481) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(2481))))  severity failure;
	assert RAM(2482) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(2482))))  severity failure;
	assert RAM(2483) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(2483))))  severity failure;
	assert RAM(2484) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(2484))))  severity failure;
	assert RAM(2485) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(2485))))  severity failure;
	assert RAM(2486) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(2486))))  severity failure;
	assert RAM(2487) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(2487))))  severity failure;
	assert RAM(2488) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(2488))))  severity failure;
	assert RAM(2489) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(2489))))  severity failure;
	assert RAM(2490) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(2490))))  severity failure;
	assert RAM(2491) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(2491))))  severity failure;
	assert RAM(2492) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(2492))))  severity failure;
	assert RAM(2493) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(2493))))  severity failure;
	assert RAM(2494) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(2494))))  severity failure;
	assert RAM(2495) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(2495))))  severity failure;
	assert RAM(2496) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(2496))))  severity failure;
	assert RAM(2497) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(2497))))  severity failure;
	assert RAM(2498) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(2498))))  severity failure;
	assert RAM(2499) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(2499))))  severity failure;
	assert RAM(2500) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(2500))))  severity failure;
	assert RAM(2501) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(2501))))  severity failure;
	assert RAM(2502) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(2502))))  severity failure;
	assert RAM(2503) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(2503))))  severity failure;
	assert RAM(2504) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(2504))))  severity failure;
	assert RAM(2505) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(2505))))  severity failure;
	assert RAM(2506) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(2506))))  severity failure;
	assert RAM(2507) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(2507))))  severity failure;
	assert RAM(2508) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(2508))))  severity failure;
	assert RAM(2509) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(2509))))  severity failure;
	assert RAM(2510) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(2510))))  severity failure;
	assert RAM(2511) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(2511))))  severity failure;
	assert RAM(2512) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(2512))))  severity failure;
	assert RAM(2513) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(2513))))  severity failure;
	assert RAM(2514) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(2514))))  severity failure;
	assert RAM(2515) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(2515))))  severity failure;
	assert RAM(2516) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(2516))))  severity failure;
	assert RAM(2517) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(2517))))  severity failure;
	assert RAM(2518) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(2518))))  severity failure;
	assert RAM(2519) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(2519))))  severity failure;
	assert RAM(2520) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(2520))))  severity failure;
	assert RAM(2521) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(2521))))  severity failure;
	assert RAM(2522) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(2522))))  severity failure;
	assert RAM(2523) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(2523))))  severity failure;
	assert RAM(2524) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(2524))))  severity failure;
	assert RAM(2525) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(2525))))  severity failure;
	assert RAM(2526) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(2526))))  severity failure;
	assert RAM(2527) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(2527))))  severity failure;
	assert RAM(2528) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(2528))))  severity failure;
	assert RAM(2529) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(2529))))  severity failure;
	assert RAM(2530) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(2530))))  severity failure;
	assert RAM(2531) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(2531))))  severity failure;
	assert RAM(2532) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(2532))))  severity failure;
	assert RAM(2533) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(2533))))  severity failure;
	assert RAM(2534) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(2534))))  severity failure;
	assert RAM(2535) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(2535))))  severity failure;
	assert RAM(2536) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(2536))))  severity failure;
	assert RAM(2537) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(2537))))  severity failure;
	assert RAM(2538) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(2538))))  severity failure;
	assert RAM(2539) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(2539))))  severity failure;
	assert RAM(2540) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(2540))))  severity failure;
	assert RAM(2541) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(2541))))  severity failure;
	assert RAM(2542) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(2542))))  severity failure;
	assert RAM(2543) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(2543))))  severity failure;
	assert RAM(2544) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(2544))))  severity failure;
	assert RAM(2545) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(2545))))  severity failure;
	assert RAM(2546) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(2546))))  severity failure;
	assert RAM(2547) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(2547))))  severity failure;
	assert RAM(2548) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(2548))))  severity failure;
	assert RAM(2549) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(2549))))  severity failure;
	assert RAM(2550) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(2550))))  severity failure;
	assert RAM(2551) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(2551))))  severity failure;
	assert RAM(2552) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(2552))))  severity failure;
	assert RAM(2553) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(2553))))  severity failure;
	assert RAM(2554) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(2554))))  severity failure;
	assert RAM(2555) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(2555))))  severity failure;
	assert RAM(2556) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(2556))))  severity failure;
	assert RAM(2557) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(2557))))  severity failure;
	assert RAM(2558) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(2558))))  severity failure;
	assert RAM(2559) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(2559))))  severity failure;
	assert RAM(2560) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(2560))))  severity failure;
	assert RAM(2561) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(2561))))  severity failure;
	assert RAM(2562) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(2562))))  severity failure;
	assert RAM(2563) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(2563))))  severity failure;
	assert RAM(2564) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(2564))))  severity failure;
	assert RAM(2565) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(2565))))  severity failure;
	assert RAM(2566) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(2566))))  severity failure;
	assert RAM(2567) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(2567))))  severity failure;
	assert RAM(2568) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(2568))))  severity failure;
	assert RAM(2569) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(2569))))  severity failure;
	assert RAM(2570) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(2570))))  severity failure;
	assert RAM(2571) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(2571))))  severity failure;
	assert RAM(2572) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(2572))))  severity failure;
	assert RAM(2573) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(2573))))  severity failure;
	assert RAM(2574) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(2574))))  severity failure;
	assert RAM(2575) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(2575))))  severity failure;
	assert RAM(2576) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(2576))))  severity failure;
	assert RAM(2577) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(2577))))  severity failure;
	assert RAM(2578) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(2578))))  severity failure;
	assert RAM(2579) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(2579))))  severity failure;
	assert RAM(2580) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(2580))))  severity failure;
	assert RAM(2581) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(2581))))  severity failure;
	assert RAM(2582) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(2582))))  severity failure;
	assert RAM(2583) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(2583))))  severity failure;
	assert RAM(2584) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(2584))))  severity failure;
	assert RAM(2585) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(2585))))  severity failure;
	assert RAM(2586) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(2586))))  severity failure;
	assert RAM(2587) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(2587))))  severity failure;
	assert RAM(2588) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(2588))))  severity failure;
	assert RAM(2589) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(2589))))  severity failure;
	assert RAM(2590) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(2590))))  severity failure;
	assert RAM(2591) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(2591))))  severity failure;
	assert RAM(2592) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(2592))))  severity failure;
	assert RAM(2593) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(2593))))  severity failure;
	assert RAM(2594) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(2594))))  severity failure;
	assert RAM(2595) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(2595))))  severity failure;
	assert RAM(2596) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(2596))))  severity failure;
	assert RAM(2597) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(2597))))  severity failure;
	assert RAM(2598) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(2598))))  severity failure;
	assert RAM(2599) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(2599))))  severity failure;
	assert RAM(2600) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(2600))))  severity failure;
	assert RAM(2601) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(2601))))  severity failure;
	assert RAM(2602) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(2602))))  severity failure;
	assert RAM(2603) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(2603))))  severity failure;
	assert RAM(2604) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(2604))))  severity failure;
	assert RAM(2605) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(2605))))  severity failure;
	assert RAM(2606) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(2606))))  severity failure;
	assert RAM(2607) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(2607))))  severity failure;
	assert RAM(2608) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(2608))))  severity failure;
	assert RAM(2609) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(2609))))  severity failure;
	assert RAM(2610) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(2610))))  severity failure;
	assert RAM(2611) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(2611))))  severity failure;
	assert RAM(2612) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(2612))))  severity failure;
	assert RAM(2613) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(2613))))  severity failure;
	assert RAM(2614) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(2614))))  severity failure;
	assert RAM(2615) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(2615))))  severity failure;
	assert RAM(2616) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(2616))))  severity failure;
	assert RAM(2617) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(2617))))  severity failure;
	assert RAM(2618) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(2618))))  severity failure;
	assert RAM(2619) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(2619))))  severity failure;
	assert RAM(2620) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(2620))))  severity failure;
	assert RAM(2621) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(2621))))  severity failure;
	assert RAM(2622) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(2622))))  severity failure;
	assert RAM(2623) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(2623))))  severity failure;
	assert RAM(2624) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(2624))))  severity failure;
	assert RAM(2625) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(2625))))  severity failure;
	assert RAM(2626) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(2626))))  severity failure;
	assert RAM(2627) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(2627))))  severity failure;
	assert RAM(2628) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(2628))))  severity failure;
	assert RAM(2629) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(2629))))  severity failure;
	assert RAM(2630) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(2630))))  severity failure;
	assert RAM(2631) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(2631))))  severity failure;
	assert RAM(2632) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(2632))))  severity failure;
	assert RAM(2633) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(2633))))  severity failure;
	assert RAM(2634) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(2634))))  severity failure;
	assert RAM(2635) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(2635))))  severity failure;
	assert RAM(2636) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(2636))))  severity failure;
	assert RAM(2637) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(2637))))  severity failure;
	assert RAM(2638) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(2638))))  severity failure;
	assert RAM(2639) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(2639))))  severity failure;
	assert RAM(2640) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(2640))))  severity failure;
	assert RAM(2641) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(2641))))  severity failure;
	assert RAM(2642) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(2642))))  severity failure;
	assert RAM(2643) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(2643))))  severity failure;
	assert RAM(2644) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(2644))))  severity failure;
	assert RAM(2645) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(2645))))  severity failure;
	assert RAM(2646) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(2646))))  severity failure;
	assert RAM(2647) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(2647))))  severity failure;
	assert RAM(2648) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(2648))))  severity failure;
	assert RAM(2649) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(2649))))  severity failure;
	assert RAM(2650) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(2650))))  severity failure;
	assert RAM(2651) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(2651))))  severity failure;
	assert RAM(2652) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(2652))))  severity failure;
	assert RAM(2653) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(2653))))  severity failure;
	assert RAM(2654) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(2654))))  severity failure;
	assert RAM(2655) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(2655))))  severity failure;
	assert RAM(2656) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(2656))))  severity failure;
	assert RAM(2657) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(2657))))  severity failure;
	assert RAM(2658) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(2658))))  severity failure;
	assert RAM(2659) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(2659))))  severity failure;
	assert RAM(2660) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(2660))))  severity failure;
	assert RAM(2661) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(2661))))  severity failure;
	assert RAM(2662) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(2662))))  severity failure;
	assert RAM(2663) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(2663))))  severity failure;
	assert RAM(2664) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(2664))))  severity failure;
	assert RAM(2665) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(2665))))  severity failure;
	assert RAM(2666) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(2666))))  severity failure;
	assert RAM(2667) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(2667))))  severity failure;
	assert RAM(2668) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(2668))))  severity failure;
	assert RAM(2669) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(2669))))  severity failure;
	assert RAM(2670) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(2670))))  severity failure;
	assert RAM(2671) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(2671))))  severity failure;
	assert RAM(2672) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(2672))))  severity failure;
	assert RAM(2673) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(2673))))  severity failure;
	assert RAM(2674) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(2674))))  severity failure;
	assert RAM(2675) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(2675))))  severity failure;
	assert RAM(2676) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(2676))))  severity failure;
	assert RAM(2677) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(2677))))  severity failure;
	assert RAM(2678) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(2678))))  severity failure;
	assert RAM(2679) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(2679))))  severity failure;
	assert RAM(2680) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(2680))))  severity failure;
	assert RAM(2681) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(2681))))  severity failure;
	assert RAM(2682) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(2682))))  severity failure;
	assert RAM(2683) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(2683))))  severity failure;
	assert RAM(2684) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(2684))))  severity failure;
	assert RAM(2685) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(2685))))  severity failure;
	assert RAM(2686) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(2686))))  severity failure;
	assert RAM(2687) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(2687))))  severity failure;
	assert RAM(2688) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(2688))))  severity failure;
	assert RAM(2689) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(2689))))  severity failure;
	assert RAM(2690) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(2690))))  severity failure;
	assert RAM(2691) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(2691))))  severity failure;
	assert RAM(2692) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(2692))))  severity failure;
	assert RAM(2693) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(2693))))  severity failure;
	assert RAM(2694) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(2694))))  severity failure;
	assert RAM(2695) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(2695))))  severity failure;
	assert RAM(2696) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(2696))))  severity failure;
	assert RAM(2697) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(2697))))  severity failure;
	assert RAM(2698) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(2698))))  severity failure;
	assert RAM(2699) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(2699))))  severity failure;
	assert RAM(2700) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(2700))))  severity failure;
	assert RAM(2701) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(2701))))  severity failure;
	assert RAM(2702) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(2702))))  severity failure;
	assert RAM(2703) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(2703))))  severity failure;
	assert RAM(2704) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(2704))))  severity failure;
	assert RAM(2705) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(2705))))  severity failure;
	assert RAM(2706) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(2706))))  severity failure;
	assert RAM(2707) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(2707))))  severity failure;
	assert RAM(2708) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(2708))))  severity failure;
	assert RAM(2709) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(2709))))  severity failure;
	assert RAM(2710) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(2710))))  severity failure;
	assert RAM(2711) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(2711))))  severity failure;
	assert RAM(2712) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(2712))))  severity failure;
	assert RAM(2713) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(2713))))  severity failure;
	assert RAM(2714) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(2714))))  severity failure;
	assert RAM(2715) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(2715))))  severity failure;
	assert RAM(2716) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(2716))))  severity failure;
	assert RAM(2717) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(2717))))  severity failure;
	assert RAM(2718) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(2718))))  severity failure;
	assert RAM(2719) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(2719))))  severity failure;
	assert RAM(2720) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(2720))))  severity failure;
	assert RAM(2721) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(2721))))  severity failure;
	assert RAM(2722) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(2722))))  severity failure;
	assert RAM(2723) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(2723))))  severity failure;
	assert RAM(2724) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(2724))))  severity failure;
	assert RAM(2725) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(2725))))  severity failure;
	assert RAM(2726) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(2726))))  severity failure;
	assert RAM(2727) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(2727))))  severity failure;
	assert RAM(2728) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(2728))))  severity failure;
	assert RAM(2729) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(2729))))  severity failure;
	assert RAM(2730) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(2730))))  severity failure;
	assert RAM(2731) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(2731))))  severity failure;
	assert RAM(2732) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(2732))))  severity failure;
	assert RAM(2733) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(2733))))  severity failure;
	assert RAM(2734) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(2734))))  severity failure;
	assert RAM(2735) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(2735))))  severity failure;
	assert RAM(2736) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(2736))))  severity failure;
	assert RAM(2737) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(2737))))  severity failure;
	assert RAM(2738) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(2738))))  severity failure;
	assert RAM(2739) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(2739))))  severity failure;
	assert RAM(2740) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(2740))))  severity failure;
	assert RAM(2741) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(2741))))  severity failure;
	assert RAM(2742) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(2742))))  severity failure;
	assert RAM(2743) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(2743))))  severity failure;
	assert RAM(2744) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(2744))))  severity failure;
	assert RAM(2745) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(2745))))  severity failure;
	assert RAM(2746) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(2746))))  severity failure;
	assert RAM(2747) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(2747))))  severity failure;
	assert RAM(2748) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(2748))))  severity failure;
	assert RAM(2749) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(2749))))  severity failure;
	assert RAM(2750) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(2750))))  severity failure;
	assert RAM(2751) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(2751))))  severity failure;
	assert RAM(2752) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(2752))))  severity failure;
	assert RAM(2753) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(2753))))  severity failure;
	assert RAM(2754) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(2754))))  severity failure;
	assert RAM(2755) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(2755))))  severity failure;
	assert RAM(2756) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(2756))))  severity failure;
	assert RAM(2757) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(2757))))  severity failure;
	assert RAM(2758) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(2758))))  severity failure;
	assert RAM(2759) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(2759))))  severity failure;
	assert RAM(2760) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(2760))))  severity failure;
	assert RAM(2761) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(2761))))  severity failure;
	assert RAM(2762) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(2762))))  severity failure;
	assert RAM(2763) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(2763))))  severity failure;
	assert RAM(2764) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(2764))))  severity failure;
	assert RAM(2765) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(2765))))  severity failure;
	assert RAM(2766) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(2766))))  severity failure;
	assert RAM(2767) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(2767))))  severity failure;
	assert RAM(2768) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(2768))))  severity failure;
	assert RAM(2769) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(2769))))  severity failure;
	assert RAM(2770) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(2770))))  severity failure;
	assert RAM(2771) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(2771))))  severity failure;
	assert RAM(2772) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(2772))))  severity failure;
	assert RAM(2773) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(2773))))  severity failure;
	assert RAM(2774) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(2774))))  severity failure;
	assert RAM(2775) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(2775))))  severity failure;
	assert RAM(2776) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(2776))))  severity failure;
	assert RAM(2777) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(2777))))  severity failure;
	assert RAM(2778) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(2778))))  severity failure;
	assert RAM(2779) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(2779))))  severity failure;
	assert RAM(2780) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(2780))))  severity failure;
	assert RAM(2781) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(2781))))  severity failure;
	assert RAM(2782) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(2782))))  severity failure;
	assert RAM(2783) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(2783))))  severity failure;
	assert RAM(2784) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(2784))))  severity failure;
	assert RAM(2785) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(2785))))  severity failure;
	assert RAM(2786) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(2786))))  severity failure;
	assert RAM(2787) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(2787))))  severity failure;
	assert RAM(2788) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(2788))))  severity failure;
	assert RAM(2789) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(2789))))  severity failure;
	assert RAM(2790) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(2790))))  severity failure;
	assert RAM(2791) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(2791))))  severity failure;
	assert RAM(2792) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(2792))))  severity failure;
	assert RAM(2793) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(2793))))  severity failure;
	assert RAM(2794) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(2794))))  severity failure;
	assert RAM(2795) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(2795))))  severity failure;
	assert RAM(2796) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(2796))))  severity failure;
	assert RAM(2797) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(2797))))  severity failure;
	assert RAM(2798) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(2798))))  severity failure;
	assert RAM(2799) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(2799))))  severity failure;
	assert RAM(2800) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(2800))))  severity failure;
	assert RAM(2801) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(2801))))  severity failure;
	assert RAM(2802) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(2802))))  severity failure;
	assert RAM(2803) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(2803))))  severity failure;
	assert RAM(2804) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(2804))))  severity failure;
	assert RAM(2805) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(2805))))  severity failure;
	assert RAM(2806) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(2806))))  severity failure;
	assert RAM(2807) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(2807))))  severity failure;
	assert RAM(2808) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(2808))))  severity failure;
	assert RAM(2809) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(2809))))  severity failure;
	assert RAM(2810) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(2810))))  severity failure;
	assert RAM(2811) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(2811))))  severity failure;
	assert RAM(2812) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(2812))))  severity failure;
	assert RAM(2813) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(2813))))  severity failure;
	assert RAM(2814) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(2814))))  severity failure;
	assert RAM(2815) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(2815))))  severity failure;
	assert RAM(2816) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(2816))))  severity failure;
	assert RAM(2817) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(2817))))  severity failure;
	assert RAM(2818) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(2818))))  severity failure;
	assert RAM(2819) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(2819))))  severity failure;
	assert RAM(2820) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(2820))))  severity failure;
	assert RAM(2821) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(2821))))  severity failure;
	assert RAM(2822) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(2822))))  severity failure;
	assert RAM(2823) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(2823))))  severity failure;
	assert RAM(2824) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(2824))))  severity failure;
	assert RAM(2825) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(2825))))  severity failure;
	assert RAM(2826) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(2826))))  severity failure;
	assert RAM(2827) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(2827))))  severity failure;
	assert RAM(2828) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(2828))))  severity failure;
	assert RAM(2829) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(2829))))  severity failure;
	assert RAM(2830) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(2830))))  severity failure;
	assert RAM(2831) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(2831))))  severity failure;
	assert RAM(2832) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(2832))))  severity failure;
	assert RAM(2833) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(2833))))  severity failure;
	assert RAM(2834) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(2834))))  severity failure;
	assert RAM(2835) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(2835))))  severity failure;
	assert RAM(2836) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(2836))))  severity failure;
	assert RAM(2837) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(2837))))  severity failure;
	assert RAM(2838) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(2838))))  severity failure;
	assert RAM(2839) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(2839))))  severity failure;
	assert RAM(2840) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(2840))))  severity failure;
	assert RAM(2841) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(2841))))  severity failure;
	assert RAM(2842) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(2842))))  severity failure;
	assert RAM(2843) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(2843))))  severity failure;
	assert RAM(2844) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(2844))))  severity failure;
	assert RAM(2845) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(2845))))  severity failure;
	assert RAM(2846) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(2846))))  severity failure;
	assert RAM(2847) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(2847))))  severity failure;
	assert RAM(2848) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(2848))))  severity failure;
	assert RAM(2849) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(2849))))  severity failure;
	assert RAM(2850) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(2850))))  severity failure;
	assert RAM(2851) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(2851))))  severity failure;
	assert RAM(2852) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(2852))))  severity failure;
	assert RAM(2853) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(2853))))  severity failure;
	assert RAM(2854) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(2854))))  severity failure;
	assert RAM(2855) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(2855))))  severity failure;
	assert RAM(2856) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(2856))))  severity failure;
	assert RAM(2857) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(2857))))  severity failure;
	assert RAM(2858) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(2858))))  severity failure;
	assert RAM(2859) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(2859))))  severity failure;
	assert RAM(2860) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(2860))))  severity failure;
	assert RAM(2861) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(2861))))  severity failure;
	assert RAM(2862) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(2862))))  severity failure;
	assert RAM(2863) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(2863))))  severity failure;
	assert RAM(2864) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(2864))))  severity failure;
	assert RAM(2865) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(2865))))  severity failure;
	assert RAM(2866) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(2866))))  severity failure;
	assert RAM(2867) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(2867))))  severity failure;
	assert RAM(2868) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(2868))))  severity failure;
	assert RAM(2869) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(2869))))  severity failure;
	assert RAM(2870) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(2870))))  severity failure;
	assert RAM(2871) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(2871))))  severity failure;
	assert RAM(2872) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(2872))))  severity failure;
	assert RAM(2873) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(2873))))  severity failure;
	assert RAM(2874) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(2874))))  severity failure;
	assert RAM(2875) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(2875))))  severity failure;
	assert RAM(2876) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(2876))))  severity failure;
	assert RAM(2877) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(2877))))  severity failure;
	assert RAM(2878) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(2878))))  severity failure;
	assert RAM(2879) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(2879))))  severity failure;
	assert RAM(2880) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(2880))))  severity failure;
	assert RAM(2881) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(2881))))  severity failure;
	assert RAM(2882) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(2882))))  severity failure;
	assert RAM(2883) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(2883))))  severity failure;
	assert RAM(2884) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(2884))))  severity failure;
	assert RAM(2885) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(2885))))  severity failure;
	assert RAM(2886) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(2886))))  severity failure;
	assert RAM(2887) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(2887))))  severity failure;
	assert RAM(2888) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(2888))))  severity failure;
	assert RAM(2889) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(2889))))  severity failure;
	assert RAM(2890) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(2890))))  severity failure;
	assert RAM(2891) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(2891))))  severity failure;
	assert RAM(2892) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(2892))))  severity failure;
	assert RAM(2893) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(2893))))  severity failure;
	assert RAM(2894) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(2894))))  severity failure;
	assert RAM(2895) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(2895))))  severity failure;
	assert RAM(2896) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(2896))))  severity failure;
	assert RAM(2897) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(2897))))  severity failure;
	assert RAM(2898) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(2898))))  severity failure;
	assert RAM(2899) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(2899))))  severity failure;
	assert RAM(2900) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(2900))))  severity failure;
	assert RAM(2901) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(2901))))  severity failure;
	assert RAM(2902) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(2902))))  severity failure;
	assert RAM(2903) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(2903))))  severity failure;
	assert RAM(2904) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(2904))))  severity failure;
	assert RAM(2905) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(2905))))  severity failure;
	assert RAM(2906) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(2906))))  severity failure;
	assert RAM(2907) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(2907))))  severity failure;
	assert RAM(2908) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(2908))))  severity failure;
	assert RAM(2909) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(2909))))  severity failure;
	assert RAM(2910) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(2910))))  severity failure;
	assert RAM(2911) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(2911))))  severity failure;
	assert RAM(2912) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(2912))))  severity failure;
	assert RAM(2913) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(2913))))  severity failure;
	assert RAM(2914) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(2914))))  severity failure;
	assert RAM(2915) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(2915))))  severity failure;
	assert RAM(2916) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(2916))))  severity failure;
	assert RAM(2917) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(2917))))  severity failure;
	assert RAM(2918) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(2918))))  severity failure;
	assert RAM(2919) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(2919))))  severity failure;
	assert RAM(2920) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(2920))))  severity failure;
	assert RAM(2921) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(2921))))  severity failure;
	assert RAM(2922) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(2922))))  severity failure;
	assert RAM(2923) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(2923))))  severity failure;
	assert RAM(2924) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(2924))))  severity failure;
	assert RAM(2925) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(2925))))  severity failure;
	assert RAM(2926) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(2926))))  severity failure;
	assert RAM(2927) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(2927))))  severity failure;
	assert RAM(2928) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(2928))))  severity failure;
	assert RAM(2929) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(2929))))  severity failure;
	assert RAM(2930) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(2930))))  severity failure;
	assert RAM(2931) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(2931))))  severity failure;
	assert RAM(2932) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(2932))))  severity failure;
	assert RAM(2933) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(2933))))  severity failure;
	assert RAM(2934) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(2934))))  severity failure;
	assert RAM(2935) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(2935))))  severity failure;
	assert RAM(2936) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(2936))))  severity failure;
	assert RAM(2937) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(2937))))  severity failure;
	assert RAM(2938) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(2938))))  severity failure;
	assert RAM(2939) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(2939))))  severity failure;
	assert RAM(2940) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(2940))))  severity failure;
	assert RAM(2941) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(2941))))  severity failure;
	assert RAM(2942) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(2942))))  severity failure;
	assert RAM(2943) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(2943))))  severity failure;
	assert RAM(2944) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(2944))))  severity failure;
	assert RAM(2945) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(2945))))  severity failure;
	assert RAM(2946) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(2946))))  severity failure;
	assert RAM(2947) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(2947))))  severity failure;
	assert RAM(2948) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(2948))))  severity failure;
	assert RAM(2949) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(2949))))  severity failure;
	assert RAM(2950) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(2950))))  severity failure;
	assert RAM(2951) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(2951))))  severity failure;
	assert RAM(2952) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(2952))))  severity failure;
	assert RAM(2953) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(2953))))  severity failure;
	assert RAM(2954) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(2954))))  severity failure;
	assert RAM(2955) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(2955))))  severity failure;
	assert RAM(2956) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(2956))))  severity failure;
	assert RAM(2957) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(2957))))  severity failure;
	assert RAM(2958) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(2958))))  severity failure;
	assert RAM(2959) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(2959))))  severity failure;
	assert RAM(2960) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(2960))))  severity failure;
	assert RAM(2961) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(2961))))  severity failure;
	assert RAM(2962) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(2962))))  severity failure;
	assert RAM(2963) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(2963))))  severity failure;
	assert RAM(2964) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(2964))))  severity failure;
	assert RAM(2965) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(2965))))  severity failure;
	assert RAM(2966) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(2966))))  severity failure;
	assert RAM(2967) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(2967))))  severity failure;
	assert RAM(2968) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(2968))))  severity failure;
	assert RAM(2969) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(2969))))  severity failure;
	assert RAM(2970) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(2970))))  severity failure;
	assert RAM(2971) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(2971))))  severity failure;
	assert RAM(2972) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(2972))))  severity failure;
	assert RAM(2973) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(2973))))  severity failure;
	assert RAM(2974) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(2974))))  severity failure;
	assert RAM(2975) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(2975))))  severity failure;
	assert RAM(2976) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(2976))))  severity failure;
	assert RAM(2977) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(2977))))  severity failure;
	assert RAM(2978) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(2978))))  severity failure;
	assert RAM(2979) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(2979))))  severity failure;
	assert RAM(2980) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(2980))))  severity failure;
	assert RAM(2981) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(2981))))  severity failure;
	assert RAM(2982) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(2982))))  severity failure;
	assert RAM(2983) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(2983))))  severity failure;
	assert RAM(2984) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(2984))))  severity failure;
	assert RAM(2985) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(2985))))  severity failure;
	assert RAM(2986) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(2986))))  severity failure;
	assert RAM(2987) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(2987))))  severity failure;
	assert RAM(2988) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(2988))))  severity failure;
	assert RAM(2989) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(2989))))  severity failure;
	assert RAM(2990) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(2990))))  severity failure;
	assert RAM(2991) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(2991))))  severity failure;
	assert RAM(2992) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(2992))))  severity failure;
	assert RAM(2993) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(2993))))  severity failure;
	assert RAM(2994) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(2994))))  severity failure;
	assert RAM(2995) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(2995))))  severity failure;
	assert RAM(2996) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(2996))))  severity failure;
	assert RAM(2997) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(2997))))  severity failure;
	assert RAM(2998) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(2998))))  severity failure;
	assert RAM(2999) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(2999))))  severity failure;
	assert RAM(3000) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(3000))))  severity failure;
	assert RAM(3001) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(3001))))  severity failure;
	assert RAM(3002) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(3002))))  severity failure;
	assert RAM(3003) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(3003))))  severity failure;
	assert RAM(3004) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(3004))))  severity failure;
	assert RAM(3005) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(3005))))  severity failure;
	assert RAM(3006) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(3006))))  severity failure;
	assert RAM(3007) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(3007))))  severity failure;
	assert RAM(3008) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(3008))))  severity failure;
	assert RAM(3009) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(3009))))  severity failure;
	assert RAM(3010) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(3010))))  severity failure;
	assert RAM(3011) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(3011))))  severity failure;
	assert RAM(3012) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(3012))))  severity failure;
	assert RAM(3013) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(3013))))  severity failure;
	assert RAM(3014) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(3014))))  severity failure;
	assert RAM(3015) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(3015))))  severity failure;
	assert RAM(3016) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(3016))))  severity failure;
	assert RAM(3017) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(3017))))  severity failure;
	assert RAM(3018) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(3018))))  severity failure;
	assert RAM(3019) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(3019))))  severity failure;
	assert RAM(3020) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(3020))))  severity failure;
	assert RAM(3021) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(3021))))  severity failure;
	assert RAM(3022) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(3022))))  severity failure;
	assert RAM(3023) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(3023))))  severity failure;
	assert RAM(3024) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(3024))))  severity failure;
	assert RAM(3025) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(3025))))  severity failure;
	assert RAM(3026) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(3026))))  severity failure;
	assert RAM(3027) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(3027))))  severity failure;
	assert RAM(3028) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(3028))))  severity failure;
	assert RAM(3029) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(3029))))  severity failure;
	assert RAM(3030) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(3030))))  severity failure;
	assert RAM(3031) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(3031))))  severity failure;
	assert RAM(3032) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(3032))))  severity failure;
	assert RAM(3033) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(3033))))  severity failure;
	assert RAM(3034) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(3034))))  severity failure;
	assert RAM(3035) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(3035))))  severity failure;
	assert RAM(3036) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(3036))))  severity failure;
	assert RAM(3037) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(3037))))  severity failure;
	assert RAM(3038) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(3038))))  severity failure;
	assert RAM(3039) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(3039))))  severity failure;
	assert RAM(3040) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(3040))))  severity failure;
	assert RAM(3041) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(3041))))  severity failure;
	assert RAM(3042) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(3042))))  severity failure;
	assert RAM(3043) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(3043))))  severity failure;
	assert RAM(3044) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(3044))))  severity failure;
	assert RAM(3045) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(3045))))  severity failure;
	assert RAM(3046) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(3046))))  severity failure;
	assert RAM(3047) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(3047))))  severity failure;
	assert RAM(3048) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(3048))))  severity failure;
	assert RAM(3049) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(3049))))  severity failure;
	assert RAM(3050) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(3050))))  severity failure;
	assert RAM(3051) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(3051))))  severity failure;
	assert RAM(3052) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(3052))))  severity failure;
	assert RAM(3053) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(3053))))  severity failure;
	assert RAM(3054) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(3054))))  severity failure;
	assert RAM(3055) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(3055))))  severity failure;
	assert RAM(3056) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(3056))))  severity failure;
	assert RAM(3057) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(3057))))  severity failure;
	assert RAM(3058) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(3058))))  severity failure;
	assert RAM(3059) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(3059))))  severity failure;
	assert RAM(3060) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(3060))))  severity failure;
	assert RAM(3061) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(3061))))  severity failure;
	assert RAM(3062) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(3062))))  severity failure;
	assert RAM(3063) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(3063))))  severity failure;
	assert RAM(3064) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(3064))))  severity failure;
	assert RAM(3065) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(3065))))  severity failure;
	assert RAM(3066) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(3066))))  severity failure;
	assert RAM(3067) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(3067))))  severity failure;
	assert RAM(3068) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(3068))))  severity failure;
	assert RAM(3069) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(3069))))  severity failure;
	assert RAM(3070) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(3070))))  severity failure;
	assert RAM(3071) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(3071))))  severity failure;
	assert RAM(3072) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(3072))))  severity failure;
	assert RAM(3073) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(3073))))  severity failure;
	assert RAM(3074) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(3074))))  severity failure;
	assert RAM(3075) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(3075))))  severity failure;
	assert RAM(3076) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(3076))))  severity failure;
	assert RAM(3077) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(3077))))  severity failure;
	assert RAM(3078) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(3078))))  severity failure;
	assert RAM(3079) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(3079))))  severity failure;
	assert RAM(3080) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(3080))))  severity failure;
	assert RAM(3081) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(3081))))  severity failure;
	assert RAM(3082) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(3082))))  severity failure;
	assert RAM(3083) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(3083))))  severity failure;
	assert RAM(3084) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(3084))))  severity failure;
	assert RAM(3085) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(3085))))  severity failure;
	assert RAM(3086) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(3086))))  severity failure;
	assert RAM(3087) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(3087))))  severity failure;
	assert RAM(3088) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(3088))))  severity failure;
	assert RAM(3089) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(3089))))  severity failure;
	assert RAM(3090) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(3090))))  severity failure;
	assert RAM(3091) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(3091))))  severity failure;
	assert RAM(3092) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(3092))))  severity failure;
	assert RAM(3093) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(3093))))  severity failure;
	assert RAM(3094) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(3094))))  severity failure;
	assert RAM(3095) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(3095))))  severity failure;
	assert RAM(3096) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(3096))))  severity failure;
	assert RAM(3097) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(3097))))  severity failure;
	assert RAM(3098) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(3098))))  severity failure;
	assert RAM(3099) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(3099))))  severity failure;
	assert RAM(3100) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(3100))))  severity failure;
	assert RAM(3101) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(3101))))  severity failure;
	assert RAM(3102) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(3102))))  severity failure;
	assert RAM(3103) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(3103))))  severity failure;
	assert RAM(3104) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(3104))))  severity failure;
	assert RAM(3105) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(3105))))  severity failure;
	assert RAM(3106) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(3106))))  severity failure;
	assert RAM(3107) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(3107))))  severity failure;
	assert RAM(3108) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(3108))))  severity failure;
	assert RAM(3109) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(3109))))  severity failure;
	assert RAM(3110) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(3110))))  severity failure;
	assert RAM(3111) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(3111))))  severity failure;
	assert RAM(3112) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(3112))))  severity failure;
	assert RAM(3113) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(3113))))  severity failure;
	assert RAM(3114) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(3114))))  severity failure;
	assert RAM(3115) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(3115))))  severity failure;
	assert RAM(3116) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(3116))))  severity failure;
	assert RAM(3117) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(3117))))  severity failure;
	assert RAM(3118) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(3118))))  severity failure;
	assert RAM(3119) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(3119))))  severity failure;
	assert RAM(3120) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(3120))))  severity failure;
	assert RAM(3121) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(3121))))  severity failure;
	assert RAM(3122) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(3122))))  severity failure;
	assert RAM(3123) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(3123))))  severity failure;
	assert RAM(3124) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(3124))))  severity failure;
	assert RAM(3125) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(3125))))  severity failure;
	assert RAM(3126) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(3126))))  severity failure;
	assert RAM(3127) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(3127))))  severity failure;
	assert RAM(3128) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(3128))))  severity failure;
	assert RAM(3129) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(3129))))  severity failure;
	assert RAM(3130) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(3130))))  severity failure;
	assert RAM(3131) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(3131))))  severity failure;
	assert RAM(3132) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(3132))))  severity failure;
	assert RAM(3133) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(3133))))  severity failure;
	assert RAM(3134) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(3134))))  severity failure;
	assert RAM(3135) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(3135))))  severity failure;
	assert RAM(3136) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(3136))))  severity failure;
	assert RAM(3137) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(3137))))  severity failure;
	assert RAM(3138) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(3138))))  severity failure;
	assert RAM(3139) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(3139))))  severity failure;
	assert RAM(3140) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(3140))))  severity failure;
	assert RAM(3141) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(3141))))  severity failure;
	assert RAM(3142) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(3142))))  severity failure;
	assert RAM(3143) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(3143))))  severity failure;
	assert RAM(3144) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(3144))))  severity failure;
	assert RAM(3145) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(3145))))  severity failure;
	assert RAM(3146) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(3146))))  severity failure;
	assert RAM(3147) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(3147))))  severity failure;
	assert RAM(3148) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(3148))))  severity failure;
	assert RAM(3149) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(3149))))  severity failure;
	assert RAM(3150) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(3150))))  severity failure;
	assert RAM(3151) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(3151))))  severity failure;
	assert RAM(3152) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(3152))))  severity failure;
	assert RAM(3153) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(3153))))  severity failure;
	assert RAM(3154) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(3154))))  severity failure;
	assert RAM(3155) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(3155))))  severity failure;
	assert RAM(3156) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(3156))))  severity failure;
	assert RAM(3157) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(3157))))  severity failure;
	assert RAM(3158) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(3158))))  severity failure;
	assert RAM(3159) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(3159))))  severity failure;
	assert RAM(3160) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(3160))))  severity failure;
	assert RAM(3161) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(3161))))  severity failure;
	assert RAM(3162) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(3162))))  severity failure;
	assert RAM(3163) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(3163))))  severity failure;
	assert RAM(3164) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(3164))))  severity failure;
	assert RAM(3165) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(3165))))  severity failure;
	assert RAM(3166) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(3166))))  severity failure;
	assert RAM(3167) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(3167))))  severity failure;
	assert RAM(3168) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(3168))))  severity failure;
	assert RAM(3169) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(3169))))  severity failure;
	assert RAM(3170) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(3170))))  severity failure;
	assert RAM(3171) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(3171))))  severity failure;
	assert RAM(3172) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(3172))))  severity failure;
	assert RAM(3173) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(3173))))  severity failure;
	assert RAM(3174) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(3174))))  severity failure;
	assert RAM(3175) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(3175))))  severity failure;
	assert RAM(3176) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(3176))))  severity failure;
	assert RAM(3177) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(3177))))  severity failure;
	assert RAM(3178) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(3178))))  severity failure;
	assert RAM(3179) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(3179))))  severity failure;
	assert RAM(3180) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(3180))))  severity failure;
	assert RAM(3181) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(3181))))  severity failure;
	assert RAM(3182) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(3182))))  severity failure;
	assert RAM(3183) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(3183))))  severity failure;
	assert RAM(3184) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(3184))))  severity failure;
	assert RAM(3185) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(3185))))  severity failure;
	assert RAM(3186) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(3186))))  severity failure;
	assert RAM(3187) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(3187))))  severity failure;
	assert RAM(3188) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(3188))))  severity failure;
	assert RAM(3189) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(3189))))  severity failure;
	assert RAM(3190) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(3190))))  severity failure;
	assert RAM(3191) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(3191))))  severity failure;
	assert RAM(3192) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(3192))))  severity failure;
	assert RAM(3193) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(3193))))  severity failure;
	assert RAM(3194) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(3194))))  severity failure;
	assert RAM(3195) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(3195))))  severity failure;
	assert RAM(3196) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(3196))))  severity failure;
	assert RAM(3197) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(3197))))  severity failure;
	assert RAM(3198) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(3198))))  severity failure;
	assert RAM(3199) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(3199))))  severity failure;
	assert RAM(3200) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(3200))))  severity failure;
	assert RAM(3201) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(3201))))  severity failure;
	assert RAM(3202) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(3202))))  severity failure;
	assert RAM(3203) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(3203))))  severity failure;
	assert RAM(3204) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(3204))))  severity failure;
	assert RAM(3205) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(3205))))  severity failure;
	assert RAM(3206) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(3206))))  severity failure;
	assert RAM(3207) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(3207))))  severity failure;
	assert RAM(3208) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(3208))))  severity failure;
	assert RAM(3209) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(3209))))  severity failure;
	assert RAM(3210) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(3210))))  severity failure;
	assert RAM(3211) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(3211))))  severity failure;
	assert RAM(3212) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(3212))))  severity failure;
	assert RAM(3213) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(3213))))  severity failure;
	assert RAM(3214) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(3214))))  severity failure;
	assert RAM(3215) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(3215))))  severity failure;
	assert RAM(3216) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(3216))))  severity failure;
	assert RAM(3217) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(3217))))  severity failure;
	assert RAM(3218) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(3218))))  severity failure;
	assert RAM(3219) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(3219))))  severity failure;
	assert RAM(3220) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(3220))))  severity failure;
	assert RAM(3221) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(3221))))  severity failure;
	assert RAM(3222) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(3222))))  severity failure;
	assert RAM(3223) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(3223))))  severity failure;
	assert RAM(3224) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(3224))))  severity failure;
	assert RAM(3225) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(3225))))  severity failure;
	assert RAM(3226) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(3226))))  severity failure;
	assert RAM(3227) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(3227))))  severity failure;
	assert RAM(3228) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(3228))))  severity failure;
	assert RAM(3229) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(3229))))  severity failure;
	assert RAM(3230) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(3230))))  severity failure;
	assert RAM(3231) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(3231))))  severity failure;
	assert RAM(3232) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(3232))))  severity failure;
	assert RAM(3233) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(3233))))  severity failure;
	assert RAM(3234) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(3234))))  severity failure;
	assert RAM(3235) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(3235))))  severity failure;
	assert RAM(3236) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(3236))))  severity failure;
	assert RAM(3237) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(3237))))  severity failure;
	assert RAM(3238) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(3238))))  severity failure;
	assert RAM(3239) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(3239))))  severity failure;
	assert RAM(3240) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(3240))))  severity failure;
	assert RAM(3241) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(3241))))  severity failure;
	assert RAM(3242) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(3242))))  severity failure;
	assert RAM(3243) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(3243))))  severity failure;
	assert RAM(3244) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(3244))))  severity failure;
	assert RAM(3245) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(3245))))  severity failure;
	assert RAM(3246) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(3246))))  severity failure;
	assert RAM(3247) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(3247))))  severity failure;
	assert RAM(3248) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(3248))))  severity failure;
	assert RAM(3249) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(3249))))  severity failure;
	assert RAM(3250) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(3250))))  severity failure;
	assert RAM(3251) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(3251))))  severity failure;
	assert RAM(3252) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(3252))))  severity failure;
	assert RAM(3253) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(3253))))  severity failure;
	assert RAM(3254) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(3254))))  severity failure;
	assert RAM(3255) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(3255))))  severity failure;
	assert RAM(3256) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(3256))))  severity failure;
	assert RAM(3257) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(3257))))  severity failure;
	assert RAM(3258) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(3258))))  severity failure;
	assert RAM(3259) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(3259))))  severity failure;
	assert RAM(3260) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(3260))))  severity failure;
	assert RAM(3261) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(3261))))  severity failure;
	assert RAM(3262) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(3262))))  severity failure;
	assert RAM(3263) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(3263))))  severity failure;
	assert RAM(3264) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(3264))))  severity failure;
	assert RAM(3265) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(3265))))  severity failure;
	assert RAM(3266) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(3266))))  severity failure;
	assert RAM(3267) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(3267))))  severity failure;
	assert RAM(3268) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(3268))))  severity failure;
	assert RAM(3269) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(3269))))  severity failure;
	assert RAM(3270) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(3270))))  severity failure;
	assert RAM(3271) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(3271))))  severity failure;
	assert RAM(3272) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(3272))))  severity failure;
	assert RAM(3273) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(3273))))  severity failure;
	assert RAM(3274) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(3274))))  severity failure;
	assert RAM(3275) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(3275))))  severity failure;
	assert RAM(3276) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(3276))))  severity failure;
	assert RAM(3277) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(3277))))  severity failure;
	assert RAM(3278) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(3278))))  severity failure;
	assert RAM(3279) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(3279))))  severity failure;
	assert RAM(3280) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(3280))))  severity failure;
	assert RAM(3281) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(3281))))  severity failure;
	assert RAM(3282) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(3282))))  severity failure;
	assert RAM(3283) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(3283))))  severity failure;
	assert RAM(3284) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(3284))))  severity failure;
	assert RAM(3285) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(3285))))  severity failure;
	assert RAM(3286) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(3286))))  severity failure;
	assert RAM(3287) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(3287))))  severity failure;
	assert RAM(3288) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(3288))))  severity failure;
	assert RAM(3289) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(3289))))  severity failure;
	assert RAM(3290) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(3290))))  severity failure;
	assert RAM(3291) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(3291))))  severity failure;
	assert RAM(3292) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(3292))))  severity failure;
	assert RAM(3293) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(3293))))  severity failure;
	assert RAM(3294) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(3294))))  severity failure;
	assert RAM(3295) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(3295))))  severity failure;
	assert RAM(3296) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(3296))))  severity failure;
	assert RAM(3297) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(3297))))  severity failure;
	assert RAM(3298) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(3298))))  severity failure;
	assert RAM(3299) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(3299))))  severity failure;
	assert RAM(3300) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(3300))))  severity failure;
	assert RAM(3301) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(3301))))  severity failure;
	assert RAM(3302) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(3302))))  severity failure;
	assert RAM(3303) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(3303))))  severity failure;
	assert RAM(3304) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(3304))))  severity failure;
	assert RAM(3305) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(3305))))  severity failure;
	assert RAM(3306) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(3306))))  severity failure;
	assert RAM(3307) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(3307))))  severity failure;
	assert RAM(3308) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(3308))))  severity failure;
	assert RAM(3309) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(3309))))  severity failure;
	assert RAM(3310) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(3310))))  severity failure;
	assert RAM(3311) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(3311))))  severity failure;
	assert RAM(3312) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(3312))))  severity failure;
	assert RAM(3313) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(3313))))  severity failure;
	assert RAM(3314) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(3314))))  severity failure;
	assert RAM(3315) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(3315))))  severity failure;
	assert RAM(3316) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(3316))))  severity failure;
	assert RAM(3317) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(3317))))  severity failure;
	assert RAM(3318) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(3318))))  severity failure;
	assert RAM(3319) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(3319))))  severity failure;
	assert RAM(3320) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(3320))))  severity failure;
	assert RAM(3321) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(3321))))  severity failure;
	assert RAM(3322) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(3322))))  severity failure;
	assert RAM(3323) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(3323))))  severity failure;
	assert RAM(3324) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(3324))))  severity failure;
	assert RAM(3325) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(3325))))  severity failure;
	assert RAM(3326) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(3326))))  severity failure;
	assert RAM(3327) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(3327))))  severity failure;
	assert RAM(3328) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(3328))))  severity failure;
	assert RAM(3329) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(3329))))  severity failure;
	assert RAM(3330) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(3330))))  severity failure;
	assert RAM(3331) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(3331))))  severity failure;
	assert RAM(3332) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(3332))))  severity failure;
	assert RAM(3333) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(3333))))  severity failure;
	assert RAM(3334) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(3334))))  severity failure;
	assert RAM(3335) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(3335))))  severity failure;
	assert RAM(3336) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(3336))))  severity failure;
	assert RAM(3337) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(3337))))  severity failure;
	assert RAM(3338) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(3338))))  severity failure;
	assert RAM(3339) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(3339))))  severity failure;
	assert RAM(3340) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(3340))))  severity failure;
	assert RAM(3341) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(3341))))  severity failure;
	assert RAM(3342) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(3342))))  severity failure;
	assert RAM(3343) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(3343))))  severity failure;
	assert RAM(3344) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(3344))))  severity failure;
	assert RAM(3345) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(3345))))  severity failure;
	assert RAM(3346) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(3346))))  severity failure;
	assert RAM(3347) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(3347))))  severity failure;
	assert RAM(3348) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(3348))))  severity failure;
	assert RAM(3349) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(3349))))  severity failure;
	assert RAM(3350) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(3350))))  severity failure;
	assert RAM(3351) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(3351))))  severity failure;
	assert RAM(3352) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(3352))))  severity failure;
	assert RAM(3353) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(3353))))  severity failure;
	assert RAM(3354) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(3354))))  severity failure;
	assert RAM(3355) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(3355))))  severity failure;
	assert RAM(3356) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(3356))))  severity failure;
	assert RAM(3357) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(3357))))  severity failure;
	assert RAM(3358) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(3358))))  severity failure;
	assert RAM(3359) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(3359))))  severity failure;
	assert RAM(3360) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(3360))))  severity failure;
	assert RAM(3361) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(3361))))  severity failure;
	assert RAM(3362) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(3362))))  severity failure;
	assert RAM(3363) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(3363))))  severity failure;
	assert RAM(3364) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(3364))))  severity failure;
	assert RAM(3365) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(3365))))  severity failure;
	assert RAM(3366) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(3366))))  severity failure;
	assert RAM(3367) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(3367))))  severity failure;
	assert RAM(3368) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(3368))))  severity failure;
	assert RAM(3369) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(3369))))  severity failure;
	assert RAM(3370) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(3370))))  severity failure;
	assert RAM(3371) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(3371))))  severity failure;
	assert RAM(3372) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(3372))))  severity failure;
	assert RAM(3373) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(3373))))  severity failure;
	assert RAM(3374) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(3374))))  severity failure;
	assert RAM(3375) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(3375))))  severity failure;
	assert RAM(3376) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(3376))))  severity failure;
	assert RAM(3377) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(3377))))  severity failure;
	assert RAM(3378) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(3378))))  severity failure;
	assert RAM(3379) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(3379))))  severity failure;
	assert RAM(3380) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(3380))))  severity failure;
	assert RAM(3381) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(3381))))  severity failure;
	assert RAM(3382) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(3382))))  severity failure;
	assert RAM(3383) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(3383))))  severity failure;
	assert RAM(3384) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(3384))))  severity failure;
	assert RAM(3385) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(3385))))  severity failure;
	assert RAM(3386) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(3386))))  severity failure;
	assert RAM(3387) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(3387))))  severity failure;
	assert RAM(3388) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(3388))))  severity failure;
	assert RAM(3389) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(3389))))  severity failure;
	assert RAM(3390) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(3390))))  severity failure;
	assert RAM(3391) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(3391))))  severity failure;
	assert RAM(3392) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(3392))))  severity failure;
	assert RAM(3393) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(3393))))  severity failure;
	assert RAM(3394) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(3394))))  severity failure;
	assert RAM(3395) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(3395))))  severity failure;
	assert RAM(3396) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(3396))))  severity failure;
	assert RAM(3397) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(3397))))  severity failure;
	assert RAM(3398) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(3398))))  severity failure;
	assert RAM(3399) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(3399))))  severity failure;
	assert RAM(3400) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(3400))))  severity failure;
	assert RAM(3401) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(3401))))  severity failure;
	assert RAM(3402) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(3402))))  severity failure;
	assert RAM(3403) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(3403))))  severity failure;
	assert RAM(3404) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(3404))))  severity failure;
	assert RAM(3405) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(3405))))  severity failure;
	assert RAM(3406) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(3406))))  severity failure;
	assert RAM(3407) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(3407))))  severity failure;
	assert RAM(3408) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(3408))))  severity failure;
	assert RAM(3409) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(3409))))  severity failure;
	assert RAM(3410) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(3410))))  severity failure;
	assert RAM(3411) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(3411))))  severity failure;
	assert RAM(3412) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(3412))))  severity failure;
	assert RAM(3413) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(3413))))  severity failure;
	assert RAM(3414) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(3414))))  severity failure;
	assert RAM(3415) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(3415))))  severity failure;
	assert RAM(3416) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(3416))))  severity failure;
	assert RAM(3417) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(3417))))  severity failure;
	assert RAM(3418) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(3418))))  severity failure;
	assert RAM(3419) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(3419))))  severity failure;
	assert RAM(3420) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(3420))))  severity failure;
	assert RAM(3421) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(3421))))  severity failure;
	assert RAM(3422) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(3422))))  severity failure;
	assert RAM(3423) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(3423))))  severity failure;
	assert RAM(3424) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(3424))))  severity failure;
	assert RAM(3425) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(3425))))  severity failure;
	assert RAM(3426) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(3426))))  severity failure;
	assert RAM(3427) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(3427))))  severity failure;
	assert RAM(3428) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(3428))))  severity failure;
	assert RAM(3429) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(3429))))  severity failure;
	assert RAM(3430) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(3430))))  severity failure;
	assert RAM(3431) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(3431))))  severity failure;
	assert RAM(3432) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(3432))))  severity failure;
	assert RAM(3433) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(3433))))  severity failure;
	assert RAM(3434) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(3434))))  severity failure;
	assert RAM(3435) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(3435))))  severity failure;
	assert RAM(3436) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(3436))))  severity failure;
	assert RAM(3437) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(3437))))  severity failure;
	assert RAM(3438) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(3438))))  severity failure;
	assert RAM(3439) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(3439))))  severity failure;
	assert RAM(3440) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(3440))))  severity failure;
	assert RAM(3441) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(3441))))  severity failure;
	assert RAM(3442) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(3442))))  severity failure;
	assert RAM(3443) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(3443))))  severity failure;
	assert RAM(3444) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(3444))))  severity failure;
	assert RAM(3445) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(3445))))  severity failure;

	assert RAM1(3612) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM1(3612))))  severity failure;
	assert RAM1(3613) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM1(3613))))  severity failure;
	assert RAM1(3614) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM1(3614))))  severity failure;
	assert RAM1(3615) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM1(3615))))  severity failure;
	assert RAM1(3616) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM1(3616))))  severity failure;
	assert RAM1(3617) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM1(3617))))  severity failure;
	assert RAM1(3618) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM1(3618))))  severity failure;
	assert RAM1(3619) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM1(3619))))  severity failure;
	assert RAM1(3620) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM1(3620))))  severity failure;
	assert RAM1(3621) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM1(3621))))  severity failure;
	assert RAM1(3622) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM1(3622))))  severity failure;
	assert RAM1(3623) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM1(3623))))  severity failure;
	assert RAM1(3624) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM1(3624))))  severity failure;
	assert RAM1(3625) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM1(3625))))  severity failure;
	assert RAM1(3626) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM1(3626))))  severity failure;
	assert RAM1(3627) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM1(3627))))  severity failure;
	assert RAM1(3628) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM1(3628))))  severity failure;
	assert RAM1(3629) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM1(3629))))  severity failure;
	assert RAM1(3630) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM1(3630))))  severity failure;
	assert RAM1(3631) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM1(3631))))  severity failure;
	assert RAM1(3632) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM1(3632))))  severity failure;
	assert RAM1(3633) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM1(3633))))  severity failure;
	assert RAM1(3634) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM1(3634))))  severity failure;
	assert RAM1(3635) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM1(3635))))  severity failure;
	assert RAM1(3636) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM1(3636))))  severity failure;
	assert RAM1(3637) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM1(3637))))  severity failure;
	assert RAM1(3638) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM1(3638))))  severity failure;
	assert RAM1(3639) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM1(3639))))  severity failure;
	assert RAM1(3640) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM1(3640))))  severity failure;
	assert RAM1(3641) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM1(3641))))  severity failure;
	assert RAM1(3642) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM1(3642))))  severity failure;
	assert RAM1(3643) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM1(3643))))  severity failure;
	assert RAM1(3644) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM1(3644))))  severity failure;
	assert RAM1(3645) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM1(3645))))  severity failure;
	assert RAM1(3646) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM1(3646))))  severity failure;
	assert RAM1(3647) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM1(3647))))  severity failure;
	assert RAM1(3648) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM1(3648))))  severity failure;
	assert RAM1(3649) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM1(3649))))  severity failure;
	assert RAM1(3650) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM1(3650))))  severity failure;
	assert RAM1(3651) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM1(3651))))  severity failure;
	assert RAM1(3652) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM1(3652))))  severity failure;
	assert RAM1(3653) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM1(3653))))  severity failure;
	assert RAM1(3654) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM1(3654))))  severity failure;
	assert RAM1(3655) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM1(3655))))  severity failure;
	assert RAM1(3656) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM1(3656))))  severity failure;
	assert RAM1(3657) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM1(3657))))  severity failure;
	assert RAM1(3658) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM1(3658))))  severity failure;
	assert RAM1(3659) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM1(3659))))  severity failure;
	assert RAM1(3660) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM1(3660))))  severity failure;
	assert RAM1(3661) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM1(3661))))  severity failure;
	assert RAM1(3662) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM1(3662))))  severity failure;
	assert RAM1(3663) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM1(3663))))  severity failure;
	assert RAM1(3664) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM1(3664))))  severity failure;
	assert RAM1(3665) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM1(3665))))  severity failure;
	assert RAM1(3666) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM1(3666))))  severity failure;
	assert RAM1(3667) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM1(3667))))  severity failure;
	assert RAM1(3668) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM1(3668))))  severity failure;
	assert RAM1(3669) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM1(3669))))  severity failure;
	assert RAM1(3670) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM1(3670))))  severity failure;
	assert RAM1(3671) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM1(3671))))  severity failure;
	assert RAM1(3672) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM1(3672))))  severity failure;
	assert RAM1(3673) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM1(3673))))  severity failure;
	assert RAM1(3674) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM1(3674))))  severity failure;
	assert RAM1(3675) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM1(3675))))  severity failure;
	assert RAM1(3676) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM1(3676))))  severity failure;
	assert RAM1(3677) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM1(3677))))  severity failure;
	assert RAM1(3678) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM1(3678))))  severity failure;
	assert RAM1(3679) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM1(3679))))  severity failure;
	assert RAM1(3680) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM1(3680))))  severity failure;
	assert RAM1(3681) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM1(3681))))  severity failure;
	assert RAM1(3682) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM1(3682))))  severity failure;
	assert RAM1(3683) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM1(3683))))  severity failure;
	assert RAM1(3684) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM1(3684))))  severity failure;
	assert RAM1(3685) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM1(3685))))  severity failure;
	assert RAM1(3686) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM1(3686))))  severity failure;
	assert RAM1(3687) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM1(3687))))  severity failure;
	assert RAM1(3688) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM1(3688))))  severity failure;
	assert RAM1(3689) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM1(3689))))  severity failure;
	assert RAM1(3690) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM1(3690))))  severity failure;
	assert RAM1(3691) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM1(3691))))  severity failure;
	assert RAM1(3692) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM1(3692))))  severity failure;
	assert RAM1(3693) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM1(3693))))  severity failure;
	assert RAM1(3694) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM1(3694))))  severity failure;
	assert RAM1(3695) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM1(3695))))  severity failure;
	assert RAM1(3696) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM1(3696))))  severity failure;
	assert RAM1(3697) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM1(3697))))  severity failure;
	assert RAM1(3698) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM1(3698))))  severity failure;
	assert RAM1(3699) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM1(3699))))  severity failure;
	assert RAM1(3700) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM1(3700))))  severity failure;
	assert RAM1(3701) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM1(3701))))  severity failure;
	assert RAM1(3702) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM1(3702))))  severity failure;
	assert RAM1(3703) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM1(3703))))  severity failure;
	assert RAM1(3704) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM1(3704))))  severity failure;
	assert RAM1(3705) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM1(3705))))  severity failure;
	assert RAM1(3706) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM1(3706))))  severity failure;
	assert RAM1(3707) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM1(3707))))  severity failure;
	assert RAM1(3708) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM1(3708))))  severity failure;
	assert RAM1(3709) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM1(3709))))  severity failure;
	assert RAM1(3710) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM1(3710))))  severity failure;
	assert RAM1(3711) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM1(3711))))  severity failure;
	assert RAM1(3712) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM1(3712))))  severity failure;
	assert RAM1(3713) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM1(3713))))  severity failure;
	assert RAM1(3714) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM1(3714))))  severity failure;
	assert RAM1(3715) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM1(3715))))  severity failure;
	assert RAM1(3716) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM1(3716))))  severity failure;
	assert RAM1(3717) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM1(3717))))  severity failure;
	assert RAM1(3718) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM1(3718))))  severity failure;
	assert RAM1(3719) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM1(3719))))  severity failure;
	assert RAM1(3720) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM1(3720))))  severity failure;
	assert RAM1(3721) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM1(3721))))  severity failure;
	assert RAM1(3722) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM1(3722))))  severity failure;
	assert RAM1(3723) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM1(3723))))  severity failure;
	assert RAM1(3724) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM1(3724))))  severity failure;
	assert RAM1(3725) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM1(3725))))  severity failure;
	assert RAM1(3726) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM1(3726))))  severity failure;
	assert RAM1(3727) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM1(3727))))  severity failure;
	assert RAM1(3728) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM1(3728))))  severity failure;
	assert RAM1(3729) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM1(3729))))  severity failure;
	assert RAM1(3730) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM1(3730))))  severity failure;
	assert RAM1(3731) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM1(3731))))  severity failure;
	assert RAM1(3732) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM1(3732))))  severity failure;
	assert RAM1(3733) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM1(3733))))  severity failure;
	assert RAM1(3734) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM1(3734))))  severity failure;
	assert RAM1(3735) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM1(3735))))  severity failure;
	assert RAM1(3736) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM1(3736))))  severity failure;
	assert RAM1(3737) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM1(3737))))  severity failure;
	assert RAM1(3738) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM1(3738))))  severity failure;
	assert RAM1(3739) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM1(3739))))  severity failure;
	assert RAM1(3740) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM1(3740))))  severity failure;
	assert RAM1(3741) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM1(3741))))  severity failure;
	assert RAM1(3742) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM1(3742))))  severity failure;
	assert RAM1(3743) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM1(3743))))  severity failure;
	assert RAM1(3744) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM1(3744))))  severity failure;
	assert RAM1(3745) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM1(3745))))  severity failure;
	assert RAM1(3746) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM1(3746))))  severity failure;
	assert RAM1(3747) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM1(3747))))  severity failure;
	assert RAM1(3748) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM1(3748))))  severity failure;
	assert RAM1(3749) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM1(3749))))  severity failure;
	assert RAM1(3750) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM1(3750))))  severity failure;
	assert RAM1(3751) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM1(3751))))  severity failure;
	assert RAM1(3752) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM1(3752))))  severity failure;
	assert RAM1(3753) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM1(3753))))  severity failure;
	assert RAM1(3754) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM1(3754))))  severity failure;
	assert RAM1(3755) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM1(3755))))  severity failure;
	assert RAM1(3756) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM1(3756))))  severity failure;
	assert RAM1(3757) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM1(3757))))  severity failure;
	assert RAM1(3758) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM1(3758))))  severity failure;
	assert RAM1(3759) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM1(3759))))  severity failure;
	assert RAM1(3760) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM1(3760))))  severity failure;
	assert RAM1(3761) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM1(3761))))  severity failure;
	assert RAM1(3762) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM1(3762))))  severity failure;
	assert RAM1(3763) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM1(3763))))  severity failure;
	assert RAM1(3764) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM1(3764))))  severity failure;
	assert RAM1(3765) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM1(3765))))  severity failure;
	assert RAM1(3766) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM1(3766))))  severity failure;
	assert RAM1(3767) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM1(3767))))  severity failure;
	assert RAM1(3768) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM1(3768))))  severity failure;
	assert RAM1(3769) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM1(3769))))  severity failure;
	assert RAM1(3770) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM1(3770))))  severity failure;
	assert RAM1(3771) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM1(3771))))  severity failure;
	assert RAM1(3772) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM1(3772))))  severity failure;
	assert RAM1(3773) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM1(3773))))  severity failure;
	assert RAM1(3774) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM1(3774))))  severity failure;
	assert RAM1(3775) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM1(3775))))  severity failure;
	assert RAM1(3776) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM1(3776))))  severity failure;
	assert RAM1(3777) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM1(3777))))  severity failure;
	assert RAM1(3778) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM1(3778))))  severity failure;
	assert RAM1(3779) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM1(3779))))  severity failure;
	assert RAM1(3780) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM1(3780))))  severity failure;
	assert RAM1(3781) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM1(3781))))  severity failure;
	assert RAM1(3782) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM1(3782))))  severity failure;
	assert RAM1(3783) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM1(3783))))  severity failure;
	assert RAM1(3784) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM1(3784))))  severity failure;
	assert RAM1(3785) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM1(3785))))  severity failure;
	assert RAM1(3786) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM1(3786))))  severity failure;
	assert RAM1(3787) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM1(3787))))  severity failure;
	assert RAM1(3788) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM1(3788))))  severity failure;
	assert RAM1(3789) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM1(3789))))  severity failure;
	assert RAM1(3790) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM1(3790))))  severity failure;
	assert RAM1(3791) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM1(3791))))  severity failure;
	assert RAM1(3792) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM1(3792))))  severity failure;
	assert RAM1(3793) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM1(3793))))  severity failure;
	assert RAM1(3794) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM1(3794))))  severity failure;
	assert RAM1(3795) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM1(3795))))  severity failure;
	assert RAM1(3796) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM1(3796))))  severity failure;
	assert RAM1(3797) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM1(3797))))  severity failure;
	assert RAM1(3798) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM1(3798))))  severity failure;
	assert RAM1(3799) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM1(3799))))  severity failure;
	assert RAM1(3800) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM1(3800))))  severity failure;
	assert RAM1(3801) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM1(3801))))  severity failure;
	assert RAM1(3802) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM1(3802))))  severity failure;
	assert RAM1(3803) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM1(3803))))  severity failure;
	assert RAM1(3804) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM1(3804))))  severity failure;
	assert RAM1(3805) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM1(3805))))  severity failure;
	assert RAM1(3806) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM1(3806))))  severity failure;
	assert RAM1(3807) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM1(3807))))  severity failure;
	assert RAM1(3808) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM1(3808))))  severity failure;
	assert RAM1(3809) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM1(3809))))  severity failure;
	assert RAM1(3810) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM1(3810))))  severity failure;
	assert RAM1(3811) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM1(3811))))  severity failure;
	assert RAM1(3812) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM1(3812))))  severity failure;
	assert RAM1(3813) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM1(3813))))  severity failure;
	assert RAM1(3814) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM1(3814))))  severity failure;
	assert RAM1(3815) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM1(3815))))  severity failure;
	assert RAM1(3816) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM1(3816))))  severity failure;
	assert RAM1(3817) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM1(3817))))  severity failure;
	assert RAM1(3818) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM1(3818))))  severity failure;
	assert RAM1(3819) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM1(3819))))  severity failure;
	assert RAM1(3820) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM1(3820))))  severity failure;
	assert RAM1(3821) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM1(3821))))  severity failure;
	assert RAM1(3822) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM1(3822))))  severity failure;
	assert RAM1(3823) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM1(3823))))  severity failure;
	assert RAM1(3824) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM1(3824))))  severity failure;
	assert RAM1(3825) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM1(3825))))  severity failure;
	assert RAM1(3826) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM1(3826))))  severity failure;
	assert RAM1(3827) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM1(3827))))  severity failure;
	assert RAM1(3828) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM1(3828))))  severity failure;
	assert RAM1(3829) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM1(3829))))  severity failure;
	assert RAM1(3830) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM1(3830))))  severity failure;
	assert RAM1(3831) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM1(3831))))  severity failure;
	assert RAM1(3832) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM1(3832))))  severity failure;
	assert RAM1(3833) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM1(3833))))  severity failure;
	assert RAM1(3834) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM1(3834))))  severity failure;
	assert RAM1(3835) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM1(3835))))  severity failure;
	assert RAM1(3836) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM1(3836))))  severity failure;
	assert RAM1(3837) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM1(3837))))  severity failure;
	assert RAM1(3838) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM1(3838))))  severity failure;
	assert RAM1(3839) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM1(3839))))  severity failure;
	assert RAM1(3840) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM1(3840))))  severity failure;
	assert RAM1(3841) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM1(3841))))  severity failure;
	assert RAM1(3842) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM1(3842))))  severity failure;
	assert RAM1(3843) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM1(3843))))  severity failure;
	assert RAM1(3844) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM1(3844))))  severity failure;
	assert RAM1(3845) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM1(3845))))  severity failure;
	assert RAM1(3846) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM1(3846))))  severity failure;
	assert RAM1(3847) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM1(3847))))  severity failure;
	assert RAM1(3848) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM1(3848))))  severity failure;
	assert RAM1(3849) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM1(3849))))  severity failure;
	assert RAM1(3850) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM1(3850))))  severity failure;
	assert RAM1(3851) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM1(3851))))  severity failure;
	assert RAM1(3852) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM1(3852))))  severity failure;
	assert RAM1(3853) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM1(3853))))  severity failure;
	assert RAM1(3854) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM1(3854))))  severity failure;
	assert RAM1(3855) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM1(3855))))  severity failure;
	assert RAM1(3856) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM1(3856))))  severity failure;
	assert RAM1(3857) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM1(3857))))  severity failure;
	assert RAM1(3858) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM1(3858))))  severity failure;
	assert RAM1(3859) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM1(3859))))  severity failure;
	assert RAM1(3860) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM1(3860))))  severity failure;
	assert RAM1(3861) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM1(3861))))  severity failure;
	assert RAM1(3862) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM1(3862))))  severity failure;
	assert RAM1(3863) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM1(3863))))  severity failure;
	assert RAM1(3864) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM1(3864))))  severity failure;
	assert RAM1(3865) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM1(3865))))  severity failure;
	assert RAM1(3866) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM1(3866))))  severity failure;
	assert RAM1(3867) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM1(3867))))  severity failure;
	assert RAM1(3868) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM1(3868))))  severity failure;
	assert RAM1(3869) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM1(3869))))  severity failure;
	assert RAM1(3870) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM1(3870))))  severity failure;
	assert RAM1(3871) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM1(3871))))  severity failure;
	assert RAM1(3872) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM1(3872))))  severity failure;
	assert RAM1(3873) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM1(3873))))  severity failure;
	assert RAM1(3874) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM1(3874))))  severity failure;
	assert RAM1(3875) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM1(3875))))  severity failure;
	assert RAM1(3876) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM1(3876))))  severity failure;
	assert RAM1(3877) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM1(3877))))  severity failure;
	assert RAM1(3878) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM1(3878))))  severity failure;
	assert RAM1(3879) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM1(3879))))  severity failure;
	assert RAM1(3880) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM1(3880))))  severity failure;
	assert RAM1(3881) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM1(3881))))  severity failure;
	assert RAM1(3882) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM1(3882))))  severity failure;
	assert RAM1(3883) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM1(3883))))  severity failure;
	assert RAM1(3884) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM1(3884))))  severity failure;
	assert RAM1(3885) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM1(3885))))  severity failure;
	assert RAM1(3886) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM1(3886))))  severity failure;
	assert RAM1(3887) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM1(3887))))  severity failure;
	assert RAM1(3888) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM1(3888))))  severity failure;
	assert RAM1(3889) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM1(3889))))  severity failure;
	assert RAM1(3890) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM1(3890))))  severity failure;
	assert RAM1(3891) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM1(3891))))  severity failure;
	assert RAM1(3892) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM1(3892))))  severity failure;
	assert RAM1(3893) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM1(3893))))  severity failure;
	assert RAM1(3894) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM1(3894))))  severity failure;
	assert RAM1(3895) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM1(3895))))  severity failure;
	assert RAM1(3896) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM1(3896))))  severity failure;
	assert RAM1(3897) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM1(3897))))  severity failure;
	assert RAM1(3898) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM1(3898))))  severity failure;
	assert RAM1(3899) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM1(3899))))  severity failure;
	assert RAM1(3900) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM1(3900))))  severity failure;
	assert RAM1(3901) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM1(3901))))  severity failure;
	assert RAM1(3902) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM1(3902))))  severity failure;
	assert RAM1(3903) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM1(3903))))  severity failure;
	assert RAM1(3904) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM1(3904))))  severity failure;
	assert RAM1(3905) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM1(3905))))  severity failure;
	assert RAM1(3906) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM1(3906))))  severity failure;
	assert RAM1(3907) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM1(3907))))  severity failure;
	assert RAM1(3908) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM1(3908))))  severity failure;
	assert RAM1(3909) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM1(3909))))  severity failure;
	assert RAM1(3910) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM1(3910))))  severity failure;
	assert RAM1(3911) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM1(3911))))  severity failure;
	assert RAM1(3912) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM1(3912))))  severity failure;
	assert RAM1(3913) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM1(3913))))  severity failure;
	assert RAM1(3914) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM1(3914))))  severity failure;
	assert RAM1(3915) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM1(3915))))  severity failure;
	assert RAM1(3916) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM1(3916))))  severity failure;
	assert RAM1(3917) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM1(3917))))  severity failure;
	assert RAM1(3918) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM1(3918))))  severity failure;
	assert RAM1(3919) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM1(3919))))  severity failure;
	assert RAM1(3920) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM1(3920))))  severity failure;
	assert RAM1(3921) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM1(3921))))  severity failure;
	assert RAM1(3922) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM1(3922))))  severity failure;
	assert RAM1(3923) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM1(3923))))  severity failure;
	assert RAM1(3924) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM1(3924))))  severity failure;
	assert RAM1(3925) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM1(3925))))  severity failure;
	assert RAM1(3926) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM1(3926))))  severity failure;
	assert RAM1(3927) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM1(3927))))  severity failure;
	assert RAM1(3928) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM1(3928))))  severity failure;
	assert RAM1(3929) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM1(3929))))  severity failure;
	assert RAM1(3930) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM1(3930))))  severity failure;
	assert RAM1(3931) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM1(3931))))  severity failure;
	assert RAM1(3932) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM1(3932))))  severity failure;
	assert RAM1(3933) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM1(3933))))  severity failure;
	assert RAM1(3934) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM1(3934))))  severity failure;
	assert RAM1(3935) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM1(3935))))  severity failure;
	assert RAM1(3936) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM1(3936))))  severity failure;
	assert RAM1(3937) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM1(3937))))  severity failure;
	assert RAM1(3938) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM1(3938))))  severity failure;
	assert RAM1(3939) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM1(3939))))  severity failure;
	assert RAM1(3940) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM1(3940))))  severity failure;
	assert RAM1(3941) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM1(3941))))  severity failure;
	assert RAM1(3942) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM1(3942))))  severity failure;
	assert RAM1(3943) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM1(3943))))  severity failure;
	assert RAM1(3944) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM1(3944))))  severity failure;
	assert RAM1(3945) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM1(3945))))  severity failure;
	assert RAM1(3946) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM1(3946))))  severity failure;
	assert RAM1(3947) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM1(3947))))  severity failure;
	assert RAM1(3948) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM1(3948))))  severity failure;
	assert RAM1(3949) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM1(3949))))  severity failure;
	assert RAM1(3950) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM1(3950))))  severity failure;
	assert RAM1(3951) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM1(3951))))  severity failure;
	assert RAM1(3952) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM1(3952))))  severity failure;
	assert RAM1(3953) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM1(3953))))  severity failure;
	assert RAM1(3954) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM1(3954))))  severity failure;
	assert RAM1(3955) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM1(3955))))  severity failure;
	assert RAM1(3956) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM1(3956))))  severity failure;
	assert RAM1(3957) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM1(3957))))  severity failure;
	assert RAM1(3958) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM1(3958))))  severity failure;
	assert RAM1(3959) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM1(3959))))  severity failure;
	assert RAM1(3960) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM1(3960))))  severity failure;
	assert RAM1(3961) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM1(3961))))  severity failure;
	assert RAM1(3962) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM1(3962))))  severity failure;
	assert RAM1(3963) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM1(3963))))  severity failure;
	assert RAM1(3964) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM1(3964))))  severity failure;
	assert RAM1(3965) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM1(3965))))  severity failure;
	assert RAM1(3966) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM1(3966))))  severity failure;
	assert RAM1(3967) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM1(3967))))  severity failure;
	assert RAM1(3968) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM1(3968))))  severity failure;
	assert RAM1(3969) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM1(3969))))  severity failure;
	assert RAM1(3970) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM1(3970))))  severity failure;
	assert RAM1(3971) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM1(3971))))  severity failure;
	assert RAM1(3972) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM1(3972))))  severity failure;
	assert RAM1(3973) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM1(3973))))  severity failure;
	assert RAM1(3974) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM1(3974))))  severity failure;
	assert RAM1(3975) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM1(3975))))  severity failure;
	assert RAM1(3976) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM1(3976))))  severity failure;
	assert RAM1(3977) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM1(3977))))  severity failure;
	assert RAM1(3978) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM1(3978))))  severity failure;
	assert RAM1(3979) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM1(3979))))  severity failure;
	assert RAM1(3980) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM1(3980))))  severity failure;
	assert RAM1(3981) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM1(3981))))  severity failure;
	assert RAM1(3982) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM1(3982))))  severity failure;
	assert RAM1(3983) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM1(3983))))  severity failure;
	assert RAM1(3984) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM1(3984))))  severity failure;
	assert RAM1(3985) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM1(3985))))  severity failure;
	assert RAM1(3986) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM1(3986))))  severity failure;
	assert RAM1(3987) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM1(3987))))  severity failure;
	assert RAM1(3988) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM1(3988))))  severity failure;
	assert RAM1(3989) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM1(3989))))  severity failure;
	assert RAM1(3990) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM1(3990))))  severity failure;
	assert RAM1(3991) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM1(3991))))  severity failure;
	assert RAM1(3992) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM1(3992))))  severity failure;
	assert RAM1(3993) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM1(3993))))  severity failure;
	assert RAM1(3994) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM1(3994))))  severity failure;
	assert RAM1(3995) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM1(3995))))  severity failure;
	assert RAM1(3996) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM1(3996))))  severity failure;
	assert RAM1(3997) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM1(3997))))  severity failure;
	assert RAM1(3998) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM1(3998))))  severity failure;
	assert RAM1(3999) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM1(3999))))  severity failure;
	assert RAM1(4000) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM1(4000))))  severity failure;
	assert RAM1(4001) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM1(4001))))  severity failure;
	assert RAM1(4002) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM1(4002))))  severity failure;
	assert RAM1(4003) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM1(4003))))  severity failure;
	assert RAM1(4004) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM1(4004))))  severity failure;
	assert RAM1(4005) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM1(4005))))  severity failure;
	assert RAM1(4006) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM1(4006))))  severity failure;
	assert RAM1(4007) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM1(4007))))  severity failure;
	assert RAM1(4008) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM1(4008))))  severity failure;
	assert RAM1(4009) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM1(4009))))  severity failure;
	assert RAM1(4010) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM1(4010))))  severity failure;
	assert RAM1(4011) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM1(4011))))  severity failure;
	assert RAM1(4012) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM1(4012))))  severity failure;
	assert RAM1(4013) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM1(4013))))  severity failure;
	assert RAM1(4014) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM1(4014))))  severity failure;
	assert RAM1(4015) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM1(4015))))  severity failure;
	assert RAM1(4016) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM1(4016))))  severity failure;
	assert RAM1(4017) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM1(4017))))  severity failure;
	assert RAM1(4018) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM1(4018))))  severity failure;
	assert RAM1(4019) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM1(4019))))  severity failure;
	assert RAM1(4020) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM1(4020))))  severity failure;
	assert RAM1(4021) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM1(4021))))  severity failure;
	assert RAM1(4022) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM1(4022))))  severity failure;
	assert RAM1(4023) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM1(4023))))  severity failure;
	assert RAM1(4024) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM1(4024))))  severity failure;
	assert RAM1(4025) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM1(4025))))  severity failure;
	assert RAM1(4026) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM1(4026))))  severity failure;
	assert RAM1(4027) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM1(4027))))  severity failure;
	assert RAM1(4028) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM1(4028))))  severity failure;
	assert RAM1(4029) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM1(4029))))  severity failure;
	assert RAM1(4030) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM1(4030))))  severity failure;
	assert RAM1(4031) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM1(4031))))  severity failure;
	assert RAM1(4032) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM1(4032))))  severity failure;
	assert RAM1(4033) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM1(4033))))  severity failure;
	assert RAM1(4034) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM1(4034))))  severity failure;
	assert RAM1(4035) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM1(4035))))  severity failure;
	assert RAM1(4036) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM1(4036))))  severity failure;
	assert RAM1(4037) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM1(4037))))  severity failure;
	assert RAM1(4038) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM1(4038))))  severity failure;
	assert RAM1(4039) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM1(4039))))  severity failure;
	assert RAM1(4040) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM1(4040))))  severity failure;
	assert RAM1(4041) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM1(4041))))  severity failure;
	assert RAM1(4042) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM1(4042))))  severity failure;
	assert RAM1(4043) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM1(4043))))  severity failure;
	assert RAM1(4044) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM1(4044))))  severity failure;
	assert RAM1(4045) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM1(4045))))  severity failure;
	assert RAM1(4046) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM1(4046))))  severity failure;
	assert RAM1(4047) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM1(4047))))  severity failure;
	assert RAM1(4048) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM1(4048))))  severity failure;
	assert RAM1(4049) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM1(4049))))  severity failure;
	assert RAM1(4050) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM1(4050))))  severity failure;
	assert RAM1(4051) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM1(4051))))  severity failure;
	assert RAM1(4052) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM1(4052))))  severity failure;
	assert RAM1(4053) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM1(4053))))  severity failure;
	assert RAM1(4054) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM1(4054))))  severity failure;
	assert RAM1(4055) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM1(4055))))  severity failure;
	assert RAM1(4056) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM1(4056))))  severity failure;
	assert RAM1(4057) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM1(4057))))  severity failure;
	assert RAM1(4058) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM1(4058))))  severity failure;
	assert RAM1(4059) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM1(4059))))  severity failure;
	assert RAM1(4060) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM1(4060))))  severity failure;
	assert RAM1(4061) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM1(4061))))  severity failure;
	assert RAM1(4062) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM1(4062))))  severity failure;
	assert RAM1(4063) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM1(4063))))  severity failure;
	assert RAM1(4064) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM1(4064))))  severity failure;
	assert RAM1(4065) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM1(4065))))  severity failure;
	assert RAM1(4066) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM1(4066))))  severity failure;
	assert RAM1(4067) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM1(4067))))  severity failure;
	assert RAM1(4068) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM1(4068))))  severity failure;
	assert RAM1(4069) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM1(4069))))  severity failure;
	assert RAM1(4070) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM1(4070))))  severity failure;
	assert RAM1(4071) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM1(4071))))  severity failure;
	assert RAM1(4072) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM1(4072))))  severity failure;
	assert RAM1(4073) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM1(4073))))  severity failure;
	assert RAM1(4074) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM1(4074))))  severity failure;
	assert RAM1(4075) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM1(4075))))  severity failure;
	assert RAM1(4076) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM1(4076))))  severity failure;
	assert RAM1(4077) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM1(4077))))  severity failure;
	assert RAM1(4078) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM1(4078))))  severity failure;
	assert RAM1(4079) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM1(4079))))  severity failure;
	assert RAM1(4080) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM1(4080))))  severity failure;
	assert RAM1(4081) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM1(4081))))  severity failure;
	assert RAM1(4082) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM1(4082))))  severity failure;
	assert RAM1(4083) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM1(4083))))  severity failure;
	assert RAM1(4084) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM1(4084))))  severity failure;
	assert RAM1(4085) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM1(4085))))  severity failure;
	assert RAM1(4086) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM1(4086))))  severity failure;
	assert RAM1(4087) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM1(4087))))  severity failure;
	assert RAM1(4088) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM1(4088))))  severity failure;
	assert RAM1(4089) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM1(4089))))  severity failure;
	assert RAM1(4090) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM1(4090))))  severity failure;
	assert RAM1(4091) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM1(4091))))  severity failure;
	assert RAM1(4092) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM1(4092))))  severity failure;
	assert RAM1(4093) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM1(4093))))  severity failure;
	assert RAM1(4094) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM1(4094))))  severity failure;
	assert RAM1(4095) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM1(4095))))  severity failure;
	assert RAM1(4096) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM1(4096))))  severity failure;
	assert RAM1(4097) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM1(4097))))  severity failure;
	assert RAM1(4098) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM1(4098))))  severity failure;
	assert RAM1(4099) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM1(4099))))  severity failure;
	assert RAM1(4100) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM1(4100))))  severity failure;
	assert RAM1(4101) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM1(4101))))  severity failure;
	assert RAM1(4102) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM1(4102))))  severity failure;
	assert RAM1(4103) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM1(4103))))  severity failure;
	assert RAM1(4104) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM1(4104))))  severity failure;
	assert RAM1(4105) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM1(4105))))  severity failure;
	assert RAM1(4106) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM1(4106))))  severity failure;
	assert RAM1(4107) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM1(4107))))  severity failure;
	assert RAM1(4108) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM1(4108))))  severity failure;
	assert RAM1(4109) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM1(4109))))  severity failure;
	assert RAM1(4110) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM1(4110))))  severity failure;
	assert RAM1(4111) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM1(4111))))  severity failure;
	assert RAM1(4112) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM1(4112))))  severity failure;
	assert RAM1(4113) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM1(4113))))  severity failure;
	assert RAM1(4114) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM1(4114))))  severity failure;
	assert RAM1(4115) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM1(4115))))  severity failure;
	assert RAM1(4116) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM1(4116))))  severity failure;
	assert RAM1(4117) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM1(4117))))  severity failure;
	assert RAM1(4118) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM1(4118))))  severity failure;
	assert RAM1(4119) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM1(4119))))  severity failure;
	assert RAM1(4120) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM1(4120))))  severity failure;
	assert RAM1(4121) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM1(4121))))  severity failure;
	assert RAM1(4122) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM1(4122))))  severity failure;
	assert RAM1(4123) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM1(4123))))  severity failure;
	assert RAM1(4124) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM1(4124))))  severity failure;
	assert RAM1(4125) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM1(4125))))  severity failure;
	assert RAM1(4126) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM1(4126))))  severity failure;
	assert RAM1(4127) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM1(4127))))  severity failure;
	assert RAM1(4128) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM1(4128))))  severity failure;
	assert RAM1(4129) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM1(4129))))  severity failure;
	assert RAM1(4130) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM1(4130))))  severity failure;
	assert RAM1(4131) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM1(4131))))  severity failure;
	assert RAM1(4132) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM1(4132))))  severity failure;
	assert RAM1(4133) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM1(4133))))  severity failure;
	assert RAM1(4134) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM1(4134))))  severity failure;
	assert RAM1(4135) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM1(4135))))  severity failure;
	assert RAM1(4136) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM1(4136))))  severity failure;
	assert RAM1(4137) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM1(4137))))  severity failure;
	assert RAM1(4138) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM1(4138))))  severity failure;
	assert RAM1(4139) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM1(4139))))  severity failure;
	assert RAM1(4140) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM1(4140))))  severity failure;
	assert RAM1(4141) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM1(4141))))  severity failure;
	assert RAM1(4142) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM1(4142))))  severity failure;
	assert RAM1(4143) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM1(4143))))  severity failure;
	assert RAM1(4144) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM1(4144))))  severity failure;
	assert RAM1(4145) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM1(4145))))  severity failure;
	assert RAM1(4146) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM1(4146))))  severity failure;
	assert RAM1(4147) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM1(4147))))  severity failure;
	assert RAM1(4148) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM1(4148))))  severity failure;
	assert RAM1(4149) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM1(4149))))  severity failure;
	assert RAM1(4150) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM1(4150))))  severity failure;
	assert RAM1(4151) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM1(4151))))  severity failure;
	assert RAM1(4152) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM1(4152))))  severity failure;
	assert RAM1(4153) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM1(4153))))  severity failure;
	assert RAM1(4154) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM1(4154))))  severity failure;
	assert RAM1(4155) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM1(4155))))  severity failure;
	assert RAM1(4156) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM1(4156))))  severity failure;
	assert RAM1(4157) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM1(4157))))  severity failure;
	assert RAM1(4158) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM1(4158))))  severity failure;
	assert RAM1(4159) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM1(4159))))  severity failure;
	assert RAM1(4160) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM1(4160))))  severity failure;
	assert RAM1(4161) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM1(4161))))  severity failure;
	assert RAM1(4162) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM1(4162))))  severity failure;
	assert RAM1(4163) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM1(4163))))  severity failure;
	assert RAM1(4164) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM1(4164))))  severity failure;
	assert RAM1(4165) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM1(4165))))  severity failure;
	assert RAM1(4166) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM1(4166))))  severity failure;
	assert RAM1(4167) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM1(4167))))  severity failure;
	assert RAM1(4168) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM1(4168))))  severity failure;
	assert RAM1(4169) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM1(4169))))  severity failure;
	assert RAM1(4170) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM1(4170))))  severity failure;
	assert RAM1(4171) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM1(4171))))  severity failure;
	assert RAM1(4172) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM1(4172))))  severity failure;
	assert RAM1(4173) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM1(4173))))  severity failure;
	assert RAM1(4174) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM1(4174))))  severity failure;
	assert RAM1(4175) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM1(4175))))  severity failure;
	assert RAM1(4176) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM1(4176))))  severity failure;
	assert RAM1(4177) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM1(4177))))  severity failure;
	assert RAM1(4178) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM1(4178))))  severity failure;
	assert RAM1(4179) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM1(4179))))  severity failure;
	assert RAM1(4180) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM1(4180))))  severity failure;
	assert RAM1(4181) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM1(4181))))  severity failure;
	assert RAM1(4182) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM1(4182))))  severity failure;
	assert RAM1(4183) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM1(4183))))  severity failure;
	assert RAM1(4184) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM1(4184))))  severity failure;
	assert RAM1(4185) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM1(4185))))  severity failure;
	assert RAM1(4186) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM1(4186))))  severity failure;
	assert RAM1(4187) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM1(4187))))  severity failure;
	assert RAM1(4188) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM1(4188))))  severity failure;
	assert RAM1(4189) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM1(4189))))  severity failure;
	assert RAM1(4190) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM1(4190))))  severity failure;
	assert RAM1(4191) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM1(4191))))  severity failure;
	assert RAM1(4192) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM1(4192))))  severity failure;
	assert RAM1(4193) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM1(4193))))  severity failure;
	assert RAM1(4194) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM1(4194))))  severity failure;
	assert RAM1(4195) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM1(4195))))  severity failure;
	assert RAM1(4196) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM1(4196))))  severity failure;
	assert RAM1(4197) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM1(4197))))  severity failure;
	assert RAM1(4198) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM1(4198))))  severity failure;
	assert RAM1(4199) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM1(4199))))  severity failure;
	assert RAM1(4200) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM1(4200))))  severity failure;
	assert RAM1(4201) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM1(4201))))  severity failure;
	assert RAM1(4202) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM1(4202))))  severity failure;
	assert RAM1(4203) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM1(4203))))  severity failure;
	assert RAM1(4204) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM1(4204))))  severity failure;
	assert RAM1(4205) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM1(4205))))  severity failure;
	assert RAM1(4206) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM1(4206))))  severity failure;
	assert RAM1(4207) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM1(4207))))  severity failure;
	assert RAM1(4208) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM1(4208))))  severity failure;
	assert RAM1(4209) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM1(4209))))  severity failure;
	assert RAM1(4210) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM1(4210))))  severity failure;
	assert RAM1(4211) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM1(4211))))  severity failure;
	assert RAM1(4212) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM1(4212))))  severity failure;
	assert RAM1(4213) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM1(4213))))  severity failure;
	assert RAM1(4214) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM1(4214))))  severity failure;
	assert RAM1(4215) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM1(4215))))  severity failure;
	assert RAM1(4216) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM1(4216))))  severity failure;
	assert RAM1(4217) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM1(4217))))  severity failure;
	assert RAM1(4218) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM1(4218))))  severity failure;
	assert RAM1(4219) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM1(4219))))  severity failure;
	assert RAM1(4220) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM1(4220))))  severity failure;
	assert RAM1(4221) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM1(4221))))  severity failure;
	assert RAM1(4222) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM1(4222))))  severity failure;
	assert RAM1(4223) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM1(4223))))  severity failure;
	assert RAM1(4224) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM1(4224))))  severity failure;
	assert RAM1(4225) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM1(4225))))  severity failure;
	assert RAM1(4226) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM1(4226))))  severity failure;
	assert RAM1(4227) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM1(4227))))  severity failure;
	assert RAM1(4228) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM1(4228))))  severity failure;
	assert RAM1(4229) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM1(4229))))  severity failure;
	assert RAM1(4230) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM1(4230))))  severity failure;
	assert RAM1(4231) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM1(4231))))  severity failure;
	assert RAM1(4232) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM1(4232))))  severity failure;
	assert RAM1(4233) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM1(4233))))  severity failure;
	assert RAM1(4234) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM1(4234))))  severity failure;
	assert RAM1(4235) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM1(4235))))  severity failure;
	assert RAM1(4236) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM1(4236))))  severity failure;
	assert RAM1(4237) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM1(4237))))  severity failure;
	assert RAM1(4238) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM1(4238))))  severity failure;
	assert RAM1(4239) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM1(4239))))  severity failure;
	assert RAM1(4240) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM1(4240))))  severity failure;
	assert RAM1(4241) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM1(4241))))  severity failure;
	assert RAM1(4242) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM1(4242))))  severity failure;
	assert RAM1(4243) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM1(4243))))  severity failure;
	assert RAM1(4244) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM1(4244))))  severity failure;
	assert RAM1(4245) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM1(4245))))  severity failure;
	assert RAM1(4246) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM1(4246))))  severity failure;
	assert RAM1(4247) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM1(4247))))  severity failure;
	assert RAM1(4248) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM1(4248))))  severity failure;
	assert RAM1(4249) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM1(4249))))  severity failure;
	assert RAM1(4250) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM1(4250))))  severity failure;
	assert RAM1(4251) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM1(4251))))  severity failure;
	assert RAM1(4252) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM1(4252))))  severity failure;
	assert RAM1(4253) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM1(4253))))  severity failure;
	assert RAM1(4254) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM1(4254))))  severity failure;
	assert RAM1(4255) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM1(4255))))  severity failure;
	assert RAM1(4256) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM1(4256))))  severity failure;
	assert RAM1(4257) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM1(4257))))  severity failure;
	assert RAM1(4258) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM1(4258))))  severity failure;
	assert RAM1(4259) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM1(4259))))  severity failure;
	assert RAM1(4260) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM1(4260))))  severity failure;
	assert RAM1(4261) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM1(4261))))  severity failure;
	assert RAM1(4262) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM1(4262))))  severity failure;
	assert RAM1(4263) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM1(4263))))  severity failure;
	assert RAM1(4264) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM1(4264))))  severity failure;
	assert RAM1(4265) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM1(4265))))  severity failure;
	assert RAM1(4266) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM1(4266))))  severity failure;
	assert RAM1(4267) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM1(4267))))  severity failure;
	assert RAM1(4268) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM1(4268))))  severity failure;
	assert RAM1(4269) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM1(4269))))  severity failure;
	assert RAM1(4270) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM1(4270))))  severity failure;
	assert RAM1(4271) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM1(4271))))  severity failure;
	assert RAM1(4272) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM1(4272))))  severity failure;
	assert RAM1(4273) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM1(4273))))  severity failure;
	assert RAM1(4274) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM1(4274))))  severity failure;
	assert RAM1(4275) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM1(4275))))  severity failure;
	assert RAM1(4276) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM1(4276))))  severity failure;
	assert RAM1(4277) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM1(4277))))  severity failure;
	assert RAM1(4278) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM1(4278))))  severity failure;
	assert RAM1(4279) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM1(4279))))  severity failure;
	assert RAM1(4280) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM1(4280))))  severity failure;
	assert RAM1(4281) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM1(4281))))  severity failure;
	assert RAM1(4282) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM1(4282))))  severity failure;
	assert RAM1(4283) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM1(4283))))  severity failure;
	assert RAM1(4284) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM1(4284))))  severity failure;
	assert RAM1(4285) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM1(4285))))  severity failure;
	assert RAM1(4286) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM1(4286))))  severity failure;
	assert RAM1(4287) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM1(4287))))  severity failure;
	assert RAM1(4288) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM1(4288))))  severity failure;
	assert RAM1(4289) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM1(4289))))  severity failure;
	assert RAM1(4290) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM1(4290))))  severity failure;
	assert RAM1(4291) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM1(4291))))  severity failure;
	assert RAM1(4292) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM1(4292))))  severity failure;
	assert RAM1(4293) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM1(4293))))  severity failure;
	assert RAM1(4294) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM1(4294))))  severity failure;
	assert RAM1(4295) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM1(4295))))  severity failure;
	assert RAM1(4296) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM1(4296))))  severity failure;
	assert RAM1(4297) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM1(4297))))  severity failure;
	assert RAM1(4298) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM1(4298))))  severity failure;
	assert RAM1(4299) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM1(4299))))  severity failure;
	assert RAM1(4300) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM1(4300))))  severity failure;
	assert RAM1(4301) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM1(4301))))  severity failure;
	assert RAM1(4302) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM1(4302))))  severity failure;
	assert RAM1(4303) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM1(4303))))  severity failure;
	assert RAM1(4304) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM1(4304))))  severity failure;
	assert RAM1(4305) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM1(4305))))  severity failure;
	assert RAM1(4306) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM1(4306))))  severity failure;
	assert RAM1(4307) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM1(4307))))  severity failure;
	assert RAM1(4308) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM1(4308))))  severity failure;
	assert RAM1(4309) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM1(4309))))  severity failure;
	assert RAM1(4310) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM1(4310))))  severity failure;
	assert RAM1(4311) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM1(4311))))  severity failure;
	assert RAM1(4312) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM1(4312))))  severity failure;
	assert RAM1(4313) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM1(4313))))  severity failure;
	assert RAM1(4314) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM1(4314))))  severity failure;
	assert RAM1(4315) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM1(4315))))  severity failure;
	assert RAM1(4316) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM1(4316))))  severity failure;
	assert RAM1(4317) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM1(4317))))  severity failure;
	assert RAM1(4318) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM1(4318))))  severity failure;
	assert RAM1(4319) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM1(4319))))  severity failure;
	assert RAM1(4320) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM1(4320))))  severity failure;
	assert RAM1(4321) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM1(4321))))  severity failure;
	assert RAM1(4322) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM1(4322))))  severity failure;
	assert RAM1(4323) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM1(4323))))  severity failure;
	assert RAM1(4324) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM1(4324))))  severity failure;
	assert RAM1(4325) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM1(4325))))  severity failure;
	assert RAM1(4326) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM1(4326))))  severity failure;
	assert RAM1(4327) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM1(4327))))  severity failure;
	assert RAM1(4328) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM1(4328))))  severity failure;
	assert RAM1(4329) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM1(4329))))  severity failure;
	assert RAM1(4330) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM1(4330))))  severity failure;
	assert RAM1(4331) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM1(4331))))  severity failure;
	assert RAM1(4332) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM1(4332))))  severity failure;
	assert RAM1(4333) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM1(4333))))  severity failure;
	assert RAM1(4334) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM1(4334))))  severity failure;
	assert RAM1(4335) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM1(4335))))  severity failure;
	assert RAM1(4336) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM1(4336))))  severity failure;
	assert RAM1(4337) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM1(4337))))  severity failure;
	assert RAM1(4338) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM1(4338))))  severity failure;
	assert RAM1(4339) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM1(4339))))  severity failure;
	assert RAM1(4340) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM1(4340))))  severity failure;
	assert RAM1(4341) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM1(4341))))  severity failure;
	assert RAM1(4342) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM1(4342))))  severity failure;
	assert RAM1(4343) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM1(4343))))  severity failure;
	assert RAM1(4344) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM1(4344))))  severity failure;
	assert RAM1(4345) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM1(4345))))  severity failure;
	assert RAM1(4346) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM1(4346))))  severity failure;
	assert RAM1(4347) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM1(4347))))  severity failure;
	assert RAM1(4348) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM1(4348))))  severity failure;
	assert RAM1(4349) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM1(4349))))  severity failure;
	assert RAM1(4350) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM1(4350))))  severity failure;
	assert RAM1(4351) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM1(4351))))  severity failure;
	assert RAM1(4352) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM1(4352))))  severity failure;
	assert RAM1(4353) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM1(4353))))  severity failure;
	assert RAM1(4354) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM1(4354))))  severity failure;
	assert RAM1(4355) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM1(4355))))  severity failure;
	assert RAM1(4356) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM1(4356))))  severity failure;
	assert RAM1(4357) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM1(4357))))  severity failure;
	assert RAM1(4358) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM1(4358))))  severity failure;
	assert RAM1(4359) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM1(4359))))  severity failure;
	assert RAM1(4360) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM1(4360))))  severity failure;
	assert RAM1(4361) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM1(4361))))  severity failure;
	assert RAM1(4362) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM1(4362))))  severity failure;
	assert RAM1(4363) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM1(4363))))  severity failure;
	assert RAM1(4364) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM1(4364))))  severity failure;
	assert RAM1(4365) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM1(4365))))  severity failure;
	assert RAM1(4366) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM1(4366))))  severity failure;
	assert RAM1(4367) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM1(4367))))  severity failure;
	assert RAM1(4368) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM1(4368))))  severity failure;
	assert RAM1(4369) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM1(4369))))  severity failure;
	assert RAM1(4370) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM1(4370))))  severity failure;
	assert RAM1(4371) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM1(4371))))  severity failure;
	assert RAM1(4372) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM1(4372))))  severity failure;
	assert RAM1(4373) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM1(4373))))  severity failure;
	assert RAM1(4374) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM1(4374))))  severity failure;
	assert RAM1(4375) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM1(4375))))  severity failure;
	assert RAM1(4376) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM1(4376))))  severity failure;
	assert RAM1(4377) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM1(4377))))  severity failure;
	assert RAM1(4378) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM1(4378))))  severity failure;
	assert RAM1(4379) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM1(4379))))  severity failure;
	assert RAM1(4380) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM1(4380))))  severity failure;
	assert RAM1(4381) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM1(4381))))  severity failure;
	assert RAM1(4382) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM1(4382))))  severity failure;
	assert RAM1(4383) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM1(4383))))  severity failure;
	assert RAM1(4384) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM1(4384))))  severity failure;
	assert RAM1(4385) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM1(4385))))  severity failure;
	assert RAM1(4386) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM1(4386))))  severity failure;
	assert RAM1(4387) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM1(4387))))  severity failure;
	assert RAM1(4388) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM1(4388))))  severity failure;
	assert RAM1(4389) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM1(4389))))  severity failure;
	assert RAM1(4390) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM1(4390))))  severity failure;
	assert RAM1(4391) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM1(4391))))  severity failure;
	assert RAM1(4392) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM1(4392))))  severity failure;
	assert RAM1(4393) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM1(4393))))  severity failure;
	assert RAM1(4394) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM1(4394))))  severity failure;
	assert RAM1(4395) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM1(4395))))  severity failure;
	assert RAM1(4396) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM1(4396))))  severity failure;
	assert RAM1(4397) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM1(4397))))  severity failure;
	assert RAM1(4398) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM1(4398))))  severity failure;
	assert RAM1(4399) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM1(4399))))  severity failure;
	assert RAM1(4400) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM1(4400))))  severity failure;
	assert RAM1(4401) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM1(4401))))  severity failure;
	assert RAM1(4402) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM1(4402))))  severity failure;
	assert RAM1(4403) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM1(4403))))  severity failure;
	assert RAM1(4404) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM1(4404))))  severity failure;
	assert RAM1(4405) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM1(4405))))  severity failure;
	assert RAM1(4406) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM1(4406))))  severity failure;
	assert RAM1(4407) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM1(4407))))  severity failure;
	assert RAM1(4408) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM1(4408))))  severity failure;
	assert RAM1(4409) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM1(4409))))  severity failure;
	assert RAM1(4410) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM1(4410))))  severity failure;
	assert RAM1(4411) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM1(4411))))  severity failure;
	assert RAM1(4412) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM1(4412))))  severity failure;
	assert RAM1(4413) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM1(4413))))  severity failure;
	assert RAM1(4414) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM1(4414))))  severity failure;
	assert RAM1(4415) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM1(4415))))  severity failure;
	assert RAM1(4416) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM1(4416))))  severity failure;
	assert RAM1(4417) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM1(4417))))  severity failure;
	assert RAM1(4418) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM1(4418))))  severity failure;
	assert RAM1(4419) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM1(4419))))  severity failure;
	assert RAM1(4420) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM1(4420))))  severity failure;
	assert RAM1(4421) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM1(4421))))  severity failure;
	assert RAM1(4422) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM1(4422))))  severity failure;
	assert RAM1(4423) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM1(4423))))  severity failure;
	assert RAM1(4424) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM1(4424))))  severity failure;
	assert RAM1(4425) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM1(4425))))  severity failure;
	assert RAM1(4426) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM1(4426))))  severity failure;
	assert RAM1(4427) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM1(4427))))  severity failure;
	assert RAM1(4428) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM1(4428))))  severity failure;
	assert RAM1(4429) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM1(4429))))  severity failure;
	assert RAM1(4430) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM1(4430))))  severity failure;
	assert RAM1(4431) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM1(4431))))  severity failure;
	assert RAM1(4432) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM1(4432))))  severity failure;
	assert RAM1(4433) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM1(4433))))  severity failure;
	assert RAM1(4434) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM1(4434))))  severity failure;
	assert RAM1(4435) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM1(4435))))  severity failure;
	assert RAM1(4436) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM1(4436))))  severity failure;
	assert RAM1(4437) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM1(4437))))  severity failure;
	assert RAM1(4438) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM1(4438))))  severity failure;
	assert RAM1(4439) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM1(4439))))  severity failure;
	assert RAM1(4440) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM1(4440))))  severity failure;
	assert RAM1(4441) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM1(4441))))  severity failure;
	assert RAM1(4442) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM1(4442))))  severity failure;
	assert RAM1(4443) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM1(4443))))  severity failure;
	assert RAM1(4444) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM1(4444))))  severity failure;
	assert RAM1(4445) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM1(4445))))  severity failure;
	assert RAM1(4446) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM1(4446))))  severity failure;
	assert RAM1(4447) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM1(4447))))  severity failure;
	assert RAM1(4448) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM1(4448))))  severity failure;
	assert RAM1(4449) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM1(4449))))  severity failure;
	assert RAM1(4450) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM1(4450))))  severity failure;
	assert RAM1(4451) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM1(4451))))  severity failure;
	assert RAM1(4452) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM1(4452))))  severity failure;
	assert RAM1(4453) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM1(4453))))  severity failure;
	assert RAM1(4454) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM1(4454))))  severity failure;
	assert RAM1(4455) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM1(4455))))  severity failure;
	assert RAM1(4456) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM1(4456))))  severity failure;
	assert RAM1(4457) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM1(4457))))  severity failure;
	assert RAM1(4458) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM1(4458))))  severity failure;
	assert RAM1(4459) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM1(4459))))  severity failure;
	assert RAM1(4460) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM1(4460))))  severity failure;
	assert RAM1(4461) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM1(4461))))  severity failure;
	assert RAM1(4462) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM1(4462))))  severity failure;
	assert RAM1(4463) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM1(4463))))  severity failure;
	assert RAM1(4464) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM1(4464))))  severity failure;
	assert RAM1(4465) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM1(4465))))  severity failure;
	assert RAM1(4466) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM1(4466))))  severity failure;
	assert RAM1(4467) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM1(4467))))  severity failure;
	assert RAM1(4468) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM1(4468))))  severity failure;
	assert RAM1(4469) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM1(4469))))  severity failure;
	assert RAM1(4470) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM1(4470))))  severity failure;
	assert RAM1(4471) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM1(4471))))  severity failure;
	assert RAM1(4472) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM1(4472))))  severity failure;
	assert RAM1(4473) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM1(4473))))  severity failure;
	assert RAM1(4474) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM1(4474))))  severity failure;
	assert RAM1(4475) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM1(4475))))  severity failure;
	assert RAM1(4476) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM1(4476))))  severity failure;
	assert RAM1(4477) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM1(4477))))  severity failure;
	assert RAM1(4478) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM1(4478))))  severity failure;
	assert RAM1(4479) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM1(4479))))  severity failure;
	assert RAM1(4480) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM1(4480))))  severity failure;
	assert RAM1(4481) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM1(4481))))  severity failure;
	assert RAM1(4482) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM1(4482))))  severity failure;
	assert RAM1(4483) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM1(4483))))  severity failure;
	assert RAM1(4484) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM1(4484))))  severity failure;
	assert RAM1(4485) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM1(4485))))  severity failure;
	assert RAM1(4486) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM1(4486))))  severity failure;
	assert RAM1(4487) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM1(4487))))  severity failure;
	assert RAM1(4488) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM1(4488))))  severity failure;
	assert RAM1(4489) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM1(4489))))  severity failure;
	assert RAM1(4490) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM1(4490))))  severity failure;
	assert RAM1(4491) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM1(4491))))  severity failure;
	assert RAM1(4492) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM1(4492))))  severity failure;
	assert RAM1(4493) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM1(4493))))  severity failure;
	assert RAM1(4494) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM1(4494))))  severity failure;
	assert RAM1(4495) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM1(4495))))  severity failure;
	assert RAM1(4496) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM1(4496))))  severity failure;
	assert RAM1(4497) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM1(4497))))  severity failure;
	assert RAM1(4498) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM1(4498))))  severity failure;
	assert RAM1(4499) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM1(4499))))  severity failure;
	assert RAM1(4500) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM1(4500))))  severity failure;
	assert RAM1(4501) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM1(4501))))  severity failure;
	assert RAM1(4502) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM1(4502))))  severity failure;
	assert RAM1(4503) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM1(4503))))  severity failure;
	assert RAM1(4504) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM1(4504))))  severity failure;
	assert RAM1(4505) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM1(4505))))  severity failure;
	assert RAM1(4506) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM1(4506))))  severity failure;
	assert RAM1(4507) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM1(4507))))  severity failure;
	assert RAM1(4508) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM1(4508))))  severity failure;
	assert RAM1(4509) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM1(4509))))  severity failure;
	assert RAM1(4510) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM1(4510))))  severity failure;
	assert RAM1(4511) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM1(4511))))  severity failure;
	assert RAM1(4512) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM1(4512))))  severity failure;
	assert RAM1(4513) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM1(4513))))  severity failure;
	assert RAM1(4514) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM1(4514))))  severity failure;
	assert RAM1(4515) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM1(4515))))  severity failure;
	assert RAM1(4516) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM1(4516))))  severity failure;
	assert RAM1(4517) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM1(4517))))  severity failure;
	assert RAM1(4518) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM1(4518))))  severity failure;
	assert RAM1(4519) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM1(4519))))  severity failure;
	assert RAM1(4520) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM1(4520))))  severity failure;
	assert RAM1(4521) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM1(4521))))  severity failure;
	assert RAM1(4522) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM1(4522))))  severity failure;
	assert RAM1(4523) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM1(4523))))  severity failure;
	assert RAM1(4524) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM1(4524))))  severity failure;
	assert RAM1(4525) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM1(4525))))  severity failure;
	assert RAM1(4526) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM1(4526))))  severity failure;
	assert RAM1(4527) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM1(4527))))  severity failure;
	assert RAM1(4528) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM1(4528))))  severity failure;
	assert RAM1(4529) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM1(4529))))  severity failure;
	assert RAM1(4530) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM1(4530))))  severity failure;
	assert RAM1(4531) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM1(4531))))  severity failure;
	assert RAM1(4532) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM1(4532))))  severity failure;
	assert RAM1(4533) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM1(4533))))  severity failure;
	assert RAM1(4534) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM1(4534))))  severity failure;
	assert RAM1(4535) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM1(4535))))  severity failure;
	assert RAM1(4536) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM1(4536))))  severity failure;
	assert RAM1(4537) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM1(4537))))  severity failure;
	assert RAM1(4538) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM1(4538))))  severity failure;
	assert RAM1(4539) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM1(4539))))  severity failure;
	assert RAM1(4540) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM1(4540))))  severity failure;
	assert RAM1(4541) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM1(4541))))  severity failure;
	assert RAM1(4542) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM1(4542))))  severity failure;
	assert RAM1(4543) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM1(4543))))  severity failure;
	assert RAM1(4544) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM1(4544))))  severity failure;
	assert RAM1(4545) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM1(4545))))  severity failure;
	assert RAM1(4546) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM1(4546))))  severity failure;
	assert RAM1(4547) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM1(4547))))  severity failure;
	assert RAM1(4548) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM1(4548))))  severity failure;
	assert RAM1(4549) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM1(4549))))  severity failure;
	assert RAM1(4550) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM1(4550))))  severity failure;
	assert RAM1(4551) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM1(4551))))  severity failure;
	assert RAM1(4552) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM1(4552))))  severity failure;
	assert RAM1(4553) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM1(4553))))  severity failure;
	assert RAM1(4554) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM1(4554))))  severity failure;
	assert RAM1(4555) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM1(4555))))  severity failure;
	assert RAM1(4556) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM1(4556))))  severity failure;
	assert RAM1(4557) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM1(4557))))  severity failure;
	assert RAM1(4558) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM1(4558))))  severity failure;
	assert RAM1(4559) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM1(4559))))  severity failure;
	assert RAM1(4560) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM1(4560))))  severity failure;
	assert RAM1(4561) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM1(4561))))  severity failure;
	assert RAM1(4562) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM1(4562))))  severity failure;
	assert RAM1(4563) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM1(4563))))  severity failure;
	assert RAM1(4564) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM1(4564))))  severity failure;
	assert RAM1(4565) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM1(4565))))  severity failure;
	assert RAM1(4566) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM1(4566))))  severity failure;
	assert RAM1(4567) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM1(4567))))  severity failure;
	assert RAM1(4568) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM1(4568))))  severity failure;
	assert RAM1(4569) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM1(4569))))  severity failure;
	assert RAM1(4570) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM1(4570))))  severity failure;
	assert RAM1(4571) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM1(4571))))  severity failure;
	assert RAM1(4572) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM1(4572))))  severity failure;
	assert RAM1(4573) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM1(4573))))  severity failure;
	assert RAM1(4574) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM1(4574))))  severity failure;
	assert RAM1(4575) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM1(4575))))  severity failure;
	assert RAM1(4576) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM1(4576))))  severity failure;
	assert RAM1(4577) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM1(4577))))  severity failure;
	assert RAM1(4578) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM1(4578))))  severity failure;
	assert RAM1(4579) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM1(4579))))  severity failure;
	assert RAM1(4580) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM1(4580))))  severity failure;
	assert RAM1(4581) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM1(4581))))  severity failure;
	assert RAM1(4582) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM1(4582))))  severity failure;
	assert RAM1(4583) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM1(4583))))  severity failure;
	assert RAM1(4584) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM1(4584))))  severity failure;
	assert RAM1(4585) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM1(4585))))  severity failure;
	assert RAM1(4586) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM1(4586))))  severity failure;
	assert RAM1(4587) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM1(4587))))  severity failure;
	assert RAM1(4588) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM1(4588))))  severity failure;
	assert RAM1(4589) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM1(4589))))  severity failure;
	assert RAM1(4590) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM1(4590))))  severity failure;
	assert RAM1(4591) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM1(4591))))  severity failure;
	assert RAM1(4592) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM1(4592))))  severity failure;
	assert RAM1(4593) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM1(4593))))  severity failure;
	assert RAM1(4594) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM1(4594))))  severity failure;
	assert RAM1(4595) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM1(4595))))  severity failure;
	assert RAM1(4596) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM1(4596))))  severity failure;
	assert RAM1(4597) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM1(4597))))  severity failure;
	assert RAM1(4598) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM1(4598))))  severity failure;
	assert RAM1(4599) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM1(4599))))  severity failure;
	assert RAM1(4600) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM1(4600))))  severity failure;
	assert RAM1(4601) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM1(4601))))  severity failure;
	assert RAM1(4602) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM1(4602))))  severity failure;
	assert RAM1(4603) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM1(4603))))  severity failure;
	assert RAM1(4604) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM1(4604))))  severity failure;
	assert RAM1(4605) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM1(4605))))  severity failure;
	assert RAM1(4606) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM1(4606))))  severity failure;
	assert RAM1(4607) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM1(4607))))  severity failure;
	assert RAM1(4608) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM1(4608))))  severity failure;
	assert RAM1(4609) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM1(4609))))  severity failure;
	assert RAM1(4610) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM1(4610))))  severity failure;
	assert RAM1(4611) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM1(4611))))  severity failure;
	assert RAM1(4612) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM1(4612))))  severity failure;
	assert RAM1(4613) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM1(4613))))  severity failure;
	assert RAM1(4614) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM1(4614))))  severity failure;
	assert RAM1(4615) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM1(4615))))  severity failure;
	assert RAM1(4616) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM1(4616))))  severity failure;
	assert RAM1(4617) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM1(4617))))  severity failure;
	assert RAM1(4618) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM1(4618))))  severity failure;
	assert RAM1(4619) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM1(4619))))  severity failure;
	assert RAM1(4620) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM1(4620))))  severity failure;
	assert RAM1(4621) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM1(4621))))  severity failure;
	assert RAM1(4622) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM1(4622))))  severity failure;
	assert RAM1(4623) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM1(4623))))  severity failure;
	assert RAM1(4624) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM1(4624))))  severity failure;
	assert RAM1(4625) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM1(4625))))  severity failure;
	assert RAM1(4626) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM1(4626))))  severity failure;
	assert RAM1(4627) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM1(4627))))  severity failure;
	assert RAM1(4628) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM1(4628))))  severity failure;
	assert RAM1(4629) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM1(4629))))  severity failure;
	assert RAM1(4630) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM1(4630))))  severity failure;
	assert RAM1(4631) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM1(4631))))  severity failure;
	assert RAM1(4632) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM1(4632))))  severity failure;
	assert RAM1(4633) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM1(4633))))  severity failure;
	assert RAM1(4634) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM1(4634))))  severity failure;
	assert RAM1(4635) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM1(4635))))  severity failure;
	assert RAM1(4636) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM1(4636))))  severity failure;
	assert RAM1(4637) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM1(4637))))  severity failure;
	assert RAM1(4638) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM1(4638))))  severity failure;
	assert RAM1(4639) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM1(4639))))  severity failure;
	assert RAM1(4640) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM1(4640))))  severity failure;
	assert RAM1(4641) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM1(4641))))  severity failure;
	assert RAM1(4642) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM1(4642))))  severity failure;
	assert RAM1(4643) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM1(4643))))  severity failure;
	assert RAM1(4644) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM1(4644))))  severity failure;
	assert RAM1(4645) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM1(4645))))  severity failure;
	assert RAM1(4646) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM1(4646))))  severity failure;
	assert RAM1(4647) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM1(4647))))  severity failure;
	assert RAM1(4648) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM1(4648))))  severity failure;
	assert RAM1(4649) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM1(4649))))  severity failure;
	assert RAM1(4650) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM1(4650))))  severity failure;
	assert RAM1(4651) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM1(4651))))  severity failure;
	assert RAM1(4652) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM1(4652))))  severity failure;
	assert RAM1(4653) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM1(4653))))  severity failure;
	assert RAM1(4654) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM1(4654))))  severity failure;
	assert RAM1(4655) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM1(4655))))  severity failure;
	assert RAM1(4656) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM1(4656))))  severity failure;
	assert RAM1(4657) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM1(4657))))  severity failure;
	assert RAM1(4658) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM1(4658))))  severity failure;
	assert RAM1(4659) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM1(4659))))  severity failure;
	assert RAM1(4660) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM1(4660))))  severity failure;
	assert RAM1(4661) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM1(4661))))  severity failure;
	assert RAM1(4662) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM1(4662))))  severity failure;
	assert RAM1(4663) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM1(4663))))  severity failure;
	assert RAM1(4664) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM1(4664))))  severity failure;
	assert RAM1(4665) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM1(4665))))  severity failure;
	assert RAM1(4666) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM1(4666))))  severity failure;
	assert RAM1(4667) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM1(4667))))  severity failure;
	assert RAM1(4668) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM1(4668))))  severity failure;
	assert RAM1(4669) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM1(4669))))  severity failure;
	assert RAM1(4670) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM1(4670))))  severity failure;
	assert RAM1(4671) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM1(4671))))  severity failure;
	assert RAM1(4672) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM1(4672))))  severity failure;
	assert RAM1(4673) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM1(4673))))  severity failure;
	assert RAM1(4674) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM1(4674))))  severity failure;
	assert RAM1(4675) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM1(4675))))  severity failure;
	assert RAM1(4676) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM1(4676))))  severity failure;
	assert RAM1(4677) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM1(4677))))  severity failure;
	assert RAM1(4678) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM1(4678))))  severity failure;
	assert RAM1(4679) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM1(4679))))  severity failure;
	assert RAM1(4680) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM1(4680))))  severity failure;
	assert RAM1(4681) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM1(4681))))  severity failure;
	assert RAM1(4682) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM1(4682))))  severity failure;
	assert RAM1(4683) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM1(4683))))  severity failure;
	assert RAM1(4684) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM1(4684))))  severity failure;
	assert RAM1(4685) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM1(4685))))  severity failure;
	assert RAM1(4686) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM1(4686))))  severity failure;
	assert RAM1(4687) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM1(4687))))  severity failure;
	assert RAM1(4688) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM1(4688))))  severity failure;
	assert RAM1(4689) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM1(4689))))  severity failure;
	assert RAM1(4690) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM1(4690))))  severity failure;
	assert RAM1(4691) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM1(4691))))  severity failure;
	assert RAM1(4692) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM1(4692))))  severity failure;
	assert RAM1(4693) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM1(4693))))  severity failure;
	assert RAM1(4694) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM1(4694))))  severity failure;
	assert RAM1(4695) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM1(4695))))  severity failure;
	assert RAM1(4696) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM1(4696))))  severity failure;
	assert RAM1(4697) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM1(4697))))  severity failure;
	assert RAM1(4698) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM1(4698))))  severity failure;
	assert RAM1(4699) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM1(4699))))  severity failure;
	assert RAM1(4700) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM1(4700))))  severity failure;
	assert RAM1(4701) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM1(4701))))  severity failure;
	assert RAM1(4702) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM1(4702))))  severity failure;
	assert RAM1(4703) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM1(4703))))  severity failure;
	assert RAM1(4704) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM1(4704))))  severity failure;
	assert RAM1(4705) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM1(4705))))  severity failure;
	assert RAM1(4706) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM1(4706))))  severity failure;
	assert RAM1(4707) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM1(4707))))  severity failure;
	assert RAM1(4708) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM1(4708))))  severity failure;
	assert RAM1(4709) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM1(4709))))  severity failure;
	assert RAM1(4710) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM1(4710))))  severity failure;
	assert RAM1(4711) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM1(4711))))  severity failure;
	assert RAM1(4712) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM1(4712))))  severity failure;
	assert RAM1(4713) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM1(4713))))  severity failure;
	assert RAM1(4714) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM1(4714))))  severity failure;
	assert RAM1(4715) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM1(4715))))  severity failure;
	assert RAM1(4716) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM1(4716))))  severity failure;
	assert RAM1(4717) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM1(4717))))  severity failure;
	assert RAM1(4718) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM1(4718))))  severity failure;
	assert RAM1(4719) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM1(4719))))  severity failure;
	assert RAM1(4720) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM1(4720))))  severity failure;
	assert RAM1(4721) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM1(4721))))  severity failure;
	assert RAM1(4722) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM1(4722))))  severity failure;
	assert RAM1(4723) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM1(4723))))  severity failure;
	assert RAM1(4724) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM1(4724))))  severity failure;
	assert RAM1(4725) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM1(4725))))  severity failure;
	assert RAM1(4726) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM1(4726))))  severity failure;
	assert RAM1(4727) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM1(4727))))  severity failure;
	assert RAM1(4728) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM1(4728))))  severity failure;
	assert RAM1(4729) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM1(4729))))  severity failure;
	assert RAM1(4730) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM1(4730))))  severity failure;
	assert RAM1(4731) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM1(4731))))  severity failure;
	assert RAM1(4732) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM1(4732))))  severity failure;
	assert RAM1(4733) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM1(4733))))  severity failure;
	assert RAM1(4734) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM1(4734))))  severity failure;
	assert RAM1(4735) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM1(4735))))  severity failure;
	assert RAM1(4736) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM1(4736))))  severity failure;
	assert RAM1(4737) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM1(4737))))  severity failure;
	assert RAM1(4738) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM1(4738))))  severity failure;
	assert RAM1(4739) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM1(4739))))  severity failure;
	assert RAM1(4740) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM1(4740))))  severity failure;
	assert RAM1(4741) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM1(4741))))  severity failure;
	assert RAM1(4742) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM1(4742))))  severity failure;
	assert RAM1(4743) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM1(4743))))  severity failure;
	assert RAM1(4744) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM1(4744))))  severity failure;
	assert RAM1(4745) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM1(4745))))  severity failure;
	assert RAM1(4746) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM1(4746))))  severity failure;
	assert RAM1(4747) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM1(4747))))  severity failure;
	assert RAM1(4748) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM1(4748))))  severity failure;
	assert RAM1(4749) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM1(4749))))  severity failure;
	assert RAM1(4750) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM1(4750))))  severity failure;
	assert RAM1(4751) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM1(4751))))  severity failure;
	assert RAM1(4752) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM1(4752))))  severity failure;
	assert RAM1(4753) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM1(4753))))  severity failure;
	assert RAM1(4754) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM1(4754))))  severity failure;
	assert RAM1(4755) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM1(4755))))  severity failure;
	assert RAM1(4756) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM1(4756))))  severity failure;
	assert RAM1(4757) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM1(4757))))  severity failure;
	assert RAM1(4758) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM1(4758))))  severity failure;
	assert RAM1(4759) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM1(4759))))  severity failure;
	assert RAM1(4760) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM1(4760))))  severity failure;
	assert RAM1(4761) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM1(4761))))  severity failure;
	assert RAM1(4762) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM1(4762))))  severity failure;
	assert RAM1(4763) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM1(4763))))  severity failure;
	assert RAM1(4764) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM1(4764))))  severity failure;
	assert RAM1(4765) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM1(4765))))  severity failure;
	assert RAM1(4766) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM1(4766))))  severity failure;
	assert RAM1(4767) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM1(4767))))  severity failure;
	assert RAM1(4768) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM1(4768))))  severity failure;
	assert RAM1(4769) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM1(4769))))  severity failure;
	assert RAM1(4770) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM1(4770))))  severity failure;
	assert RAM1(4771) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM1(4771))))  severity failure;
	assert RAM1(4772) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM1(4772))))  severity failure;
	assert RAM1(4773) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM1(4773))))  severity failure;
	assert RAM1(4774) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM1(4774))))  severity failure;
	assert RAM1(4775) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM1(4775))))  severity failure;
	assert RAM1(4776) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM1(4776))))  severity failure;
	assert RAM1(4777) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM1(4777))))  severity failure;
	assert RAM1(4778) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM1(4778))))  severity failure;
	assert RAM1(4779) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM1(4779))))  severity failure;
	assert RAM1(4780) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM1(4780))))  severity failure;
	assert RAM1(4781) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM1(4781))))  severity failure;
	assert RAM1(4782) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM1(4782))))  severity failure;
	assert RAM1(4783) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM1(4783))))  severity failure;
	assert RAM1(4784) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM1(4784))))  severity failure;
	assert RAM1(4785) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM1(4785))))  severity failure;
	assert RAM1(4786) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM1(4786))))  severity failure;
	assert RAM1(4787) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM1(4787))))  severity failure;
	assert RAM1(4788) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM1(4788))))  severity failure;
	assert RAM1(4789) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM1(4789))))  severity failure;
	assert RAM1(4790) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM1(4790))))  severity failure;
	assert RAM1(4791) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM1(4791))))  severity failure;
	assert RAM1(4792) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM1(4792))))  severity failure;
	assert RAM1(4793) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM1(4793))))  severity failure;
	assert RAM1(4794) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM1(4794))))  severity failure;
	assert RAM1(4795) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM1(4795))))  severity failure;
	assert RAM1(4796) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM1(4796))))  severity failure;
	assert RAM1(4797) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM1(4797))))  severity failure;
	assert RAM1(4798) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM1(4798))))  severity failure;
	assert RAM1(4799) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM1(4799))))  severity failure;
	assert RAM1(4800) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM1(4800))))  severity failure;
	assert RAM1(4801) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM1(4801))))  severity failure;
	assert RAM1(4802) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM1(4802))))  severity failure;
	assert RAM1(4803) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM1(4803))))  severity failure;
	assert RAM1(4804) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM1(4804))))  severity failure;
	assert RAM1(4805) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM1(4805))))  severity failure;
	assert RAM1(4806) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM1(4806))))  severity failure;
	assert RAM1(4807) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM1(4807))))  severity failure;
	assert RAM1(4808) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM1(4808))))  severity failure;
	assert RAM1(4809) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM1(4809))))  severity failure;
	assert RAM1(4810) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM1(4810))))  severity failure;
	assert RAM1(4811) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM1(4811))))  severity failure;
	assert RAM1(4812) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM1(4812))))  severity failure;
	assert RAM1(4813) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM1(4813))))  severity failure;
	assert RAM1(4814) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM1(4814))))  severity failure;
	assert RAM1(4815) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM1(4815))))  severity failure;
	assert RAM1(4816) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM1(4816))))  severity failure;
	assert RAM1(4817) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM1(4817))))  severity failure;
	assert RAM1(4818) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM1(4818))))  severity failure;
	assert RAM1(4819) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM1(4819))))  severity failure;
	assert RAM1(4820) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM1(4820))))  severity failure;
	assert RAM1(4821) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM1(4821))))  severity failure;
	assert RAM1(4822) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM1(4822))))  severity failure;
	assert RAM1(4823) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM1(4823))))  severity failure;
	assert RAM1(4824) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM1(4824))))  severity failure;
	assert RAM1(4825) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM1(4825))))  severity failure;
	assert RAM1(4826) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM1(4826))))  severity failure;
	assert RAM1(4827) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM1(4827))))  severity failure;
	assert RAM1(4828) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM1(4828))))  severity failure;
	assert RAM1(4829) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM1(4829))))  severity failure;
	assert RAM1(4830) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM1(4830))))  severity failure;
	assert RAM1(4831) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM1(4831))))  severity failure;
	assert RAM1(4832) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM1(4832))))  severity failure;
	assert RAM1(4833) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM1(4833))))  severity failure;
	assert RAM1(4834) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM1(4834))))  severity failure;
	assert RAM1(4835) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM1(4835))))  severity failure;
	assert RAM1(4836) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM1(4836))))  severity failure;
	assert RAM1(4837) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM1(4837))))  severity failure;
	assert RAM1(4838) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM1(4838))))  severity failure;
	assert RAM1(4839) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM1(4839))))  severity failure;
	assert RAM1(4840) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM1(4840))))  severity failure;
	assert RAM1(4841) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM1(4841))))  severity failure;
	assert RAM1(4842) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM1(4842))))  severity failure;
	assert RAM1(4843) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM1(4843))))  severity failure;
	assert RAM1(4844) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM1(4844))))  severity failure;
	assert RAM1(4845) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM1(4845))))  severity failure;
	assert RAM1(4846) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM1(4846))))  severity failure;
	assert RAM1(4847) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM1(4847))))  severity failure;
	assert RAM1(4848) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM1(4848))))  severity failure;
	assert RAM1(4849) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM1(4849))))  severity failure;
	assert RAM1(4850) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM1(4850))))  severity failure;
	assert RAM1(4851) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM1(4851))))  severity failure;
	assert RAM1(4852) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM1(4852))))  severity failure;
	assert RAM1(4853) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM1(4853))))  severity failure;
	assert RAM1(4854) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM1(4854))))  severity failure;
	assert RAM1(4855) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM1(4855))))  severity failure;
	assert RAM1(4856) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM1(4856))))  severity failure;
	assert RAM1(4857) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM1(4857))))  severity failure;
	assert RAM1(4858) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM1(4858))))  severity failure;
	assert RAM1(4859) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM1(4859))))  severity failure;
	assert RAM1(4860) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM1(4860))))  severity failure;
	assert RAM1(4861) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM1(4861))))  severity failure;
	assert RAM1(4862) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM1(4862))))  severity failure;
	assert RAM1(4863) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM1(4863))))  severity failure;
	assert RAM1(4864) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM1(4864))))  severity failure;
	assert RAM1(4865) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM1(4865))))  severity failure;
	assert RAM1(4866) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM1(4866))))  severity failure;
	assert RAM1(4867) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM1(4867))))  severity failure;
	assert RAM1(4868) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM1(4868))))  severity failure;
	assert RAM1(4869) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM1(4869))))  severity failure;
	assert RAM1(4870) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM1(4870))))  severity failure;
	assert RAM1(4871) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM1(4871))))  severity failure;
	assert RAM1(4872) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM1(4872))))  severity failure;
	assert RAM1(4873) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM1(4873))))  severity failure;
	assert RAM1(4874) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM1(4874))))  severity failure;
	assert RAM1(4875) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM1(4875))))  severity failure;
	assert RAM1(4876) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM1(4876))))  severity failure;
	assert RAM1(4877) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM1(4877))))  severity failure;
	assert RAM1(4878) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM1(4878))))  severity failure;
	assert RAM1(4879) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM1(4879))))  severity failure;
	assert RAM1(4880) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM1(4880))))  severity failure;
	assert RAM1(4881) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM1(4881))))  severity failure;
	assert RAM1(4882) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM1(4882))))  severity failure;
	assert RAM1(4883) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM1(4883))))  severity failure;
	assert RAM1(4884) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM1(4884))))  severity failure;
	assert RAM1(4885) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM1(4885))))  severity failure;
	assert RAM1(4886) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM1(4886))))  severity failure;
	assert RAM1(4887) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM1(4887))))  severity failure;
	assert RAM1(4888) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM1(4888))))  severity failure;
	assert RAM1(4889) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM1(4889))))  severity failure;
	assert RAM1(4890) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM1(4890))))  severity failure;
	assert RAM1(4891) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM1(4891))))  severity failure;
	assert RAM1(4892) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM1(4892))))  severity failure;
	assert RAM1(4893) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM1(4893))))  severity failure;
	assert RAM1(4894) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM1(4894))))  severity failure;
	assert RAM1(4895) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM1(4895))))  severity failure;
	assert RAM1(4896) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM1(4896))))  severity failure;
	assert RAM1(4897) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM1(4897))))  severity failure;
	assert RAM1(4898) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM1(4898))))  severity failure;
	assert RAM1(4899) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM1(4899))))  severity failure;
	assert RAM1(4900) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM1(4900))))  severity failure;
	assert RAM1(4901) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM1(4901))))  severity failure;
	assert RAM1(4902) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM1(4902))))  severity failure;
	assert RAM1(4903) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM1(4903))))  severity failure;
	assert RAM1(4904) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM1(4904))))  severity failure;
	assert RAM1(4905) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM1(4905))))  severity failure;
	assert RAM1(4906) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM1(4906))))  severity failure;
	assert RAM1(4907) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM1(4907))))  severity failure;
	assert RAM1(4908) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM1(4908))))  severity failure;
	assert RAM1(4909) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM1(4909))))  severity failure;
	assert RAM1(4910) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM1(4910))))  severity failure;
	assert RAM1(4911) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM1(4911))))  severity failure;
	assert RAM1(4912) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM1(4912))))  severity failure;
	assert RAM1(4913) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM1(4913))))  severity failure;
	assert RAM1(4914) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM1(4914))))  severity failure;
	assert RAM1(4915) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM1(4915))))  severity failure;
	assert RAM1(4916) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM1(4916))))  severity failure;
	assert RAM1(4917) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM1(4917))))  severity failure;
	assert RAM1(4918) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM1(4918))))  severity failure;
	assert RAM1(4919) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM1(4919))))  severity failure;
	assert RAM1(4920) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM1(4920))))  severity failure;
	assert RAM1(4921) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM1(4921))))  severity failure;
	assert RAM1(4922) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM1(4922))))  severity failure;
	assert RAM1(4923) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM1(4923))))  severity failure;
	assert RAM1(4924) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM1(4924))))  severity failure;
	assert RAM1(4925) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM1(4925))))  severity failure;
	assert RAM1(4926) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM1(4926))))  severity failure;
	assert RAM1(4927) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM1(4927))))  severity failure;
	assert RAM1(4928) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM1(4928))))  severity failure;
	assert RAM1(4929) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM1(4929))))  severity failure;
	assert RAM1(4930) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM1(4930))))  severity failure;
	assert RAM1(4931) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM1(4931))))  severity failure;
	assert RAM1(4932) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM1(4932))))  severity failure;
	assert RAM1(4933) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM1(4933))))  severity failure;
	assert RAM1(4934) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM1(4934))))  severity failure;
	assert RAM1(4935) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM1(4935))))  severity failure;
	assert RAM1(4936) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM1(4936))))  severity failure;
	assert RAM1(4937) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM1(4937))))  severity failure;
	assert RAM1(4938) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM1(4938))))  severity failure;
	assert RAM1(4939) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM1(4939))))  severity failure;
	assert RAM1(4940) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM1(4940))))  severity failure;
	assert RAM1(4941) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM1(4941))))  severity failure;
	assert RAM1(4942) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM1(4942))))  severity failure;
	assert RAM1(4943) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM1(4943))))  severity failure;
	assert RAM1(4944) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM1(4944))))  severity failure;
	assert RAM1(4945) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM1(4945))))  severity failure;
	assert RAM1(4946) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM1(4946))))  severity failure;
	assert RAM1(4947) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM1(4947))))  severity failure;
	assert RAM1(4948) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM1(4948))))  severity failure;
	assert RAM1(4949) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM1(4949))))  severity failure;
	assert RAM1(4950) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM1(4950))))  severity failure;
	assert RAM1(4951) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM1(4951))))  severity failure;
	assert RAM1(4952) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM1(4952))))  severity failure;
	assert RAM1(4953) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM1(4953))))  severity failure;
	assert RAM1(4954) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM1(4954))))  severity failure;
	assert RAM1(4955) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM1(4955))))  severity failure;
	assert RAM1(4956) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM1(4956))))  severity failure;
	assert RAM1(4957) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM1(4957))))  severity failure;
	assert RAM1(4958) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM1(4958))))  severity failure;
	assert RAM1(4959) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM1(4959))))  severity failure;
	assert RAM1(4960) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM1(4960))))  severity failure;
	assert RAM1(4961) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM1(4961))))  severity failure;
	assert RAM1(4962) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM1(4962))))  severity failure;
	assert RAM1(4963) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM1(4963))))  severity failure;
	assert RAM1(4964) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM1(4964))))  severity failure;
	assert RAM1(4965) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM1(4965))))  severity failure;
	assert RAM1(4966) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM1(4966))))  severity failure;
	assert RAM1(4967) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM1(4967))))  severity failure;
	assert RAM1(4968) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM1(4968))))  severity failure;
	assert RAM1(4969) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM1(4969))))  severity failure;
	assert RAM1(4970) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM1(4970))))  severity failure;
	assert RAM1(4971) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM1(4971))))  severity failure;
	assert RAM1(4972) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM1(4972))))  severity failure;
	assert RAM1(4973) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM1(4973))))  severity failure;
	assert RAM1(4974) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM1(4974))))  severity failure;
	assert RAM1(4975) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM1(4975))))  severity failure;
	assert RAM1(4976) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM1(4976))))  severity failure;
	assert RAM1(4977) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM1(4977))))  severity failure;
	assert RAM1(4978) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM1(4978))))  severity failure;
	assert RAM1(4979) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM1(4979))))  severity failure;
	assert RAM1(4980) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM1(4980))))  severity failure;
	assert RAM1(4981) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM1(4981))))  severity failure;
	assert RAM1(4982) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM1(4982))))  severity failure;
	assert RAM1(4983) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM1(4983))))  severity failure;
	assert RAM1(4984) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM1(4984))))  severity failure;
	assert RAM1(4985) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM1(4985))))  severity failure;
	assert RAM1(4986) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM1(4986))))  severity failure;
	assert RAM1(4987) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM1(4987))))  severity failure;
	assert RAM1(4988) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM1(4988))))  severity failure;
	assert RAM1(4989) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM1(4989))))  severity failure;
	assert RAM1(4990) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM1(4990))))  severity failure;
	assert RAM1(4991) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM1(4991))))  severity failure;
	assert RAM1(4992) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM1(4992))))  severity failure;
	assert RAM1(4993) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM1(4993))))  severity failure;
	assert RAM1(4994) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM1(4994))))  severity failure;
	assert RAM1(4995) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM1(4995))))  severity failure;
	assert RAM1(4996) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM1(4996))))  severity failure;
	assert RAM1(4997) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM1(4997))))  severity failure;
	assert RAM1(4998) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM1(4998))))  severity failure;
	assert RAM1(4999) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM1(4999))))  severity failure;
	assert RAM1(5000) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM1(5000))))  severity failure;
	assert RAM1(5001) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM1(5001))))  severity failure;
	assert RAM1(5002) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM1(5002))))  severity failure;
	assert RAM1(5003) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM1(5003))))  severity failure;
	assert RAM1(5004) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM1(5004))))  severity failure;
	assert RAM1(5005) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM1(5005))))  severity failure;
	assert RAM1(5006) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM1(5006))))  severity failure;
	assert RAM1(5007) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM1(5007))))  severity failure;
	assert RAM1(5008) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM1(5008))))  severity failure;
	assert RAM1(5009) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM1(5009))))  severity failure;
	assert RAM1(5010) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM1(5010))))  severity failure;
	assert RAM1(5011) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM1(5011))))  severity failure;
	assert RAM1(5012) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM1(5012))))  severity failure;
	assert RAM1(5013) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM1(5013))))  severity failure;
	assert RAM1(5014) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM1(5014))))  severity failure;
	assert RAM1(5015) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM1(5015))))  severity failure;
	assert RAM1(5016) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM1(5016))))  severity failure;
	assert RAM1(5017) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM1(5017))))  severity failure;
	assert RAM1(5018) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM1(5018))))  severity failure;
	assert RAM1(5019) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM1(5019))))  severity failure;
	assert RAM1(5020) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM1(5020))))  severity failure;
	assert RAM1(5021) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM1(5021))))  severity failure;
	assert RAM1(5022) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM1(5022))))  severity failure;
	assert RAM1(5023) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM1(5023))))  severity failure;
	assert RAM1(5024) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM1(5024))))  severity failure;
	assert RAM1(5025) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM1(5025))))  severity failure;
	assert RAM1(5026) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM1(5026))))  severity failure;
	assert RAM1(5027) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM1(5027))))  severity failure;
	assert RAM1(5028) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM1(5028))))  severity failure;
	assert RAM1(5029) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM1(5029))))  severity failure;
	assert RAM1(5030) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM1(5030))))  severity failure;
	assert RAM1(5031) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM1(5031))))  severity failure;
	assert RAM1(5032) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM1(5032))))  severity failure;
	assert RAM1(5033) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM1(5033))))  severity failure;
	assert RAM1(5034) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM1(5034))))  severity failure;
	assert RAM1(5035) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM1(5035))))  severity failure;
	assert RAM1(5036) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM1(5036))))  severity failure;
	assert RAM1(5037) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM1(5037))))  severity failure;
	assert RAM1(5038) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM1(5038))))  severity failure;
	assert RAM1(5039) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM1(5039))))  severity failure;
	assert RAM1(5040) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM1(5040))))  severity failure;
	assert RAM1(5041) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM1(5041))))  severity failure;
	assert RAM1(5042) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM1(5042))))  severity failure;
	assert RAM1(5043) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM1(5043))))  severity failure;
	assert RAM1(5044) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM1(5044))))  severity failure;
	assert RAM1(5045) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM1(5045))))  severity failure;
	assert RAM1(5046) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM1(5046))))  severity failure;
	assert RAM1(5047) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM1(5047))))  severity failure;
	assert RAM1(5048) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM1(5048))))  severity failure;
	assert RAM1(5049) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM1(5049))))  severity failure;
	assert RAM1(5050) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM1(5050))))  severity failure;
	assert RAM1(5051) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM1(5051))))  severity failure;
	assert RAM1(5052) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM1(5052))))  severity failure;
	assert RAM1(5053) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM1(5053))))  severity failure;
	assert RAM1(5054) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM1(5054))))  severity failure;
	assert RAM1(5055) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM1(5055))))  severity failure;
	assert RAM1(5056) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM1(5056))))  severity failure;
	assert RAM1(5057) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM1(5057))))  severity failure;
	assert RAM1(5058) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM1(5058))))  severity failure;
	assert RAM1(5059) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM1(5059))))  severity failure;
	assert RAM1(5060) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM1(5060))))  severity failure;
	assert RAM1(5061) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM1(5061))))  severity failure;
	assert RAM1(5062) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM1(5062))))  severity failure;
	assert RAM1(5063) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM1(5063))))  severity failure;
	assert RAM1(5064) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM1(5064))))  severity failure;
	assert RAM1(5065) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM1(5065))))  severity failure;
	assert RAM1(5066) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM1(5066))))  severity failure;
	assert RAM1(5067) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM1(5067))))  severity failure;
	assert RAM1(5068) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM1(5068))))  severity failure;
	assert RAM1(5069) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM1(5069))))  severity failure;
	assert RAM1(5070) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM1(5070))))  severity failure;
	assert RAM1(5071) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM1(5071))))  severity failure;
	assert RAM1(5072) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM1(5072))))  severity failure;
	assert RAM1(5073) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM1(5073))))  severity failure;
	assert RAM1(5074) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM1(5074))))  severity failure;
	assert RAM1(5075) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM1(5075))))  severity failure;
	assert RAM1(5076) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM1(5076))))  severity failure;
	assert RAM1(5077) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM1(5077))))  severity failure;
	assert RAM1(5078) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM1(5078))))  severity failure;
	assert RAM1(5079) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM1(5079))))  severity failure;
	assert RAM1(5080) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM1(5080))))  severity failure;
	assert RAM1(5081) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM1(5081))))  severity failure;
	assert RAM1(5082) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM1(5082))))  severity failure;
	assert RAM1(5083) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM1(5083))))  severity failure;
	assert RAM1(5084) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM1(5084))))  severity failure;
	assert RAM1(5085) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM1(5085))))  severity failure;
	assert RAM1(5086) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM1(5086))))  severity failure;
	assert RAM1(5087) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM1(5087))))  severity failure;
	assert RAM1(5088) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM1(5088))))  severity failure;
	assert RAM1(5089) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM1(5089))))  severity failure;
	assert RAM1(5090) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM1(5090))))  severity failure;
	assert RAM1(5091) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM1(5091))))  severity failure;
	assert RAM1(5092) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM1(5092))))  severity failure;
	assert RAM1(5093) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM1(5093))))  severity failure;
	assert RAM1(5094) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM1(5094))))  severity failure;
	assert RAM1(5095) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM1(5095))))  severity failure;
	assert RAM1(5096) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM1(5096))))  severity failure;
	assert RAM1(5097) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM1(5097))))  severity failure;
	assert RAM1(5098) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM1(5098))))  severity failure;
	assert RAM1(5099) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM1(5099))))  severity failure;
	assert RAM1(5100) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM1(5100))))  severity failure;
	assert RAM1(5101) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM1(5101))))  severity failure;
	assert RAM1(5102) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM1(5102))))  severity failure;
	assert RAM1(5103) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM1(5103))))  severity failure;
	assert RAM1(5104) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM1(5104))))  severity failure;
	assert RAM1(5105) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM1(5105))))  severity failure;
	assert RAM1(5106) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM1(5106))))  severity failure;
	assert RAM1(5107) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM1(5107))))  severity failure;
	assert RAM1(5108) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM1(5108))))  severity failure;
	assert RAM1(5109) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM1(5109))))  severity failure;
	assert RAM1(5110) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM1(5110))))  severity failure;
	assert RAM1(5111) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM1(5111))))  severity failure;
	assert RAM1(5112) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM1(5112))))  severity failure;
	assert RAM1(5113) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM1(5113))))  severity failure;
	assert RAM1(5114) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM1(5114))))  severity failure;
	assert RAM1(5115) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM1(5115))))  severity failure;
	assert RAM1(5116) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM1(5116))))  severity failure;
	assert RAM1(5117) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM1(5117))))  severity failure;
	assert RAM1(5118) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM1(5118))))  severity failure;
	assert RAM1(5119) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM1(5119))))  severity failure;
	assert RAM1(5120) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM1(5120))))  severity failure;
	assert RAM1(5121) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM1(5121))))  severity failure;
	assert RAM1(5122) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM1(5122))))  severity failure;
	assert RAM1(5123) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM1(5123))))  severity failure;
	assert RAM1(5124) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM1(5124))))  severity failure;
	assert RAM1(5125) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM1(5125))))  severity failure;
	assert RAM1(5126) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM1(5126))))  severity failure;
	assert RAM1(5127) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM1(5127))))  severity failure;
	assert RAM1(5128) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM1(5128))))  severity failure;
	assert RAM1(5129) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM1(5129))))  severity failure;
	assert RAM1(5130) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM1(5130))))  severity failure;
	assert RAM1(5131) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM1(5131))))  severity failure;
	assert RAM1(5132) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM1(5132))))  severity failure;
	assert RAM1(5133) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM1(5133))))  severity failure;
	assert RAM1(5134) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM1(5134))))  severity failure;
	assert RAM1(5135) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM1(5135))))  severity failure;
	assert RAM1(5136) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM1(5136))))  severity failure;
	assert RAM1(5137) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM1(5137))))  severity failure;
	assert RAM1(5138) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM1(5138))))  severity failure;
	assert RAM1(5139) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM1(5139))))  severity failure;
	assert RAM1(5140) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM1(5140))))  severity failure;
	assert RAM1(5141) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM1(5141))))  severity failure;
	assert RAM1(5142) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM1(5142))))  severity failure;
	assert RAM1(5143) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM1(5143))))  severity failure;
	assert RAM1(5144) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM1(5144))))  severity failure;
	assert RAM1(5145) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM1(5145))))  severity failure;
	assert RAM1(5146) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM1(5146))))  severity failure;
	assert RAM1(5147) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM1(5147))))  severity failure;
	assert RAM1(5148) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM1(5148))))  severity failure;
	assert RAM1(5149) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM1(5149))))  severity failure;
	assert RAM1(5150) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM1(5150))))  severity failure;
	assert RAM1(5151) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM1(5151))))  severity failure;
	assert RAM1(5152) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM1(5152))))  severity failure;
	assert RAM1(5153) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM1(5153))))  severity failure;
	assert RAM1(5154) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM1(5154))))  severity failure;
	assert RAM1(5155) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM1(5155))))  severity failure;
	assert RAM1(5156) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM1(5156))))  severity failure;
	assert RAM1(5157) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM1(5157))))  severity failure;
	assert RAM1(5158) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM1(5158))))  severity failure;
	assert RAM1(5159) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM1(5159))))  severity failure;
	assert RAM1(5160) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM1(5160))))  severity failure;
	assert RAM1(5161) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM1(5161))))  severity failure;
	assert RAM1(5162) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM1(5162))))  severity failure;
	assert RAM1(5163) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM1(5163))))  severity failure;
	assert RAM1(5164) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM1(5164))))  severity failure;
	assert RAM1(5165) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM1(5165))))  severity failure;
	assert RAM1(5166) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM1(5166))))  severity failure;
	assert RAM1(5167) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM1(5167))))  severity failure;
	assert RAM1(5168) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM1(5168))))  severity failure;
	assert RAM1(5169) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM1(5169))))  severity failure;
	assert RAM1(5170) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM1(5170))))  severity failure;
	assert RAM1(5171) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM1(5171))))  severity failure;
	assert RAM1(5172) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM1(5172))))  severity failure;
	assert RAM1(5173) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM1(5173))))  severity failure;
	assert RAM1(5174) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM1(5174))))  severity failure;
	assert RAM1(5175) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM1(5175))))  severity failure;
	assert RAM1(5176) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM1(5176))))  severity failure;
	assert RAM1(5177) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM1(5177))))  severity failure;
	assert RAM1(5178) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM1(5178))))  severity failure;
	assert RAM1(5179) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM1(5179))))  severity failure;
	assert RAM1(5180) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM1(5180))))  severity failure;
	assert RAM1(5181) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM1(5181))))  severity failure;
	assert RAM1(5182) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM1(5182))))  severity failure;
	assert RAM1(5183) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM1(5183))))  severity failure;
	assert RAM1(5184) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM1(5184))))  severity failure;
	assert RAM1(5185) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM1(5185))))  severity failure;
	assert RAM1(5186) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM1(5186))))  severity failure;
	assert RAM1(5187) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM1(5187))))  severity failure;
	assert RAM1(5188) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM1(5188))))  severity failure;
	assert RAM1(5189) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM1(5189))))  severity failure;
	assert RAM1(5190) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM1(5190))))  severity failure;
	assert RAM1(5191) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM1(5191))))  severity failure;
	assert RAM1(5192) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM1(5192))))  severity failure;
	assert RAM1(5193) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM1(5193))))  severity failure;
	assert RAM1(5194) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM1(5194))))  severity failure;
	assert RAM1(5195) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM1(5195))))  severity failure;
	assert RAM1(5196) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM1(5196))))  severity failure;
	assert RAM1(5197) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM1(5197))))  severity failure;
	assert RAM1(5198) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM1(5198))))  severity failure;
	assert RAM1(5199) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM1(5199))))  severity failure;
	assert RAM1(5200) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM1(5200))))  severity failure;
	assert RAM1(5201) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM1(5201))))  severity failure;
	assert RAM1(5202) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM1(5202))))  severity failure;
	assert RAM1(5203) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM1(5203))))  severity failure;
	assert RAM1(5204) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM1(5204))))  severity failure;
	assert RAM1(5205) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM1(5205))))  severity failure;
	assert RAM1(5206) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM1(5206))))  severity failure;
	assert RAM1(5207) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM1(5207))))  severity failure;
	assert RAM1(5208) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM1(5208))))  severity failure;
	assert RAM1(5209) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM1(5209))))  severity failure;
	assert RAM1(5210) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM1(5210))))  severity failure;
	assert RAM1(5211) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM1(5211))))  severity failure;
	assert RAM1(5212) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM1(5212))))  severity failure;
	assert RAM1(5213) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM1(5213))))  severity failure;
	assert RAM1(5214) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM1(5214))))  severity failure;
	assert RAM1(5215) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM1(5215))))  severity failure;
	assert RAM1(5216) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM1(5216))))  severity failure;
	assert RAM1(5217) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM1(5217))))  severity failure;
	assert RAM1(5218) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM1(5218))))  severity failure;
	assert RAM1(5219) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM1(5219))))  severity failure;
	assert RAM1(5220) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM1(5220))))  severity failure;
	assert RAM1(5221) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM1(5221))))  severity failure;
	assert RAM1(5222) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM1(5222))))  severity failure;
	assert RAM1(5223) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM1(5223))))  severity failure;
	assert RAM1(5224) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM1(5224))))  severity failure;
	assert RAM1(5225) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM1(5225))))  severity failure;
	assert RAM1(5226) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM1(5226))))  severity failure;
	assert RAM1(5227) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM1(5227))))  severity failure;
	assert RAM1(5228) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM1(5228))))  severity failure;
	assert RAM1(5229) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM1(5229))))  severity failure;
	assert RAM1(5230) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM1(5230))))  severity failure;
	assert RAM1(5231) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM1(5231))))  severity failure;
	assert RAM1(5232) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM1(5232))))  severity failure;
	assert RAM1(5233) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM1(5233))))  severity failure;
	assert RAM1(5234) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM1(5234))))  severity failure;
	assert RAM1(5235) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM1(5235))))  severity failure;
	assert RAM1(5236) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM1(5236))))  severity failure;
	assert RAM1(5237) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM1(5237))))  severity failure;
	assert RAM1(5238) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM1(5238))))  severity failure;
	assert RAM1(5239) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM1(5239))))  severity failure;
	assert RAM1(5240) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM1(5240))))  severity failure;
	assert RAM1(5241) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM1(5241))))  severity failure;
	assert RAM1(5242) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM1(5242))))  severity failure;
	assert RAM1(5243) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM1(5243))))  severity failure;
	assert RAM1(5244) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM1(5244))))  severity failure;
	assert RAM1(5245) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM1(5245))))  severity failure;
	assert RAM1(5246) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM1(5246))))  severity failure;
	assert RAM1(5247) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM1(5247))))  severity failure;
	assert RAM1(5248) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM1(5248))))  severity failure;
	assert RAM1(5249) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM1(5249))))  severity failure;
	assert RAM1(5250) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM1(5250))))  severity failure;
	assert RAM1(5251) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM1(5251))))  severity failure;
	assert RAM1(5252) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM1(5252))))  severity failure;
	assert RAM1(5253) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM1(5253))))  severity failure;
	assert RAM1(5254) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM1(5254))))  severity failure;
	assert RAM1(5255) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM1(5255))))  severity failure;
	assert RAM1(5256) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM1(5256))))  severity failure;
	assert RAM1(5257) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM1(5257))))  severity failure;
	assert RAM1(5258) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM1(5258))))  severity failure;
	assert RAM1(5259) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM1(5259))))  severity failure;
	assert RAM1(5260) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM1(5260))))  severity failure;
	assert RAM1(5261) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM1(5261))))  severity failure;
	assert RAM1(5262) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM1(5262))))  severity failure;
	assert RAM1(5263) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM1(5263))))  severity failure;
	assert RAM1(5264) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM1(5264))))  severity failure;
	assert RAM1(5265) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM1(5265))))  severity failure;
	assert RAM1(5266) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM1(5266))))  severity failure;
	assert RAM1(5267) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM1(5267))))  severity failure;
	assert RAM1(5268) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM1(5268))))  severity failure;
	assert RAM1(5269) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM1(5269))))  severity failure;
	assert RAM1(5270) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM1(5270))))  severity failure;
	assert RAM1(5271) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM1(5271))))  severity failure;
	assert RAM1(5272) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM1(5272))))  severity failure;
	assert RAM1(5273) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM1(5273))))  severity failure;
	assert RAM1(5274) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM1(5274))))  severity failure;
	assert RAM1(5275) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM1(5275))))  severity failure;
	assert RAM1(5276) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM1(5276))))  severity failure;
	assert RAM1(5277) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM1(5277))))  severity failure;
	assert RAM1(5278) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM1(5278))))  severity failure;
	assert RAM1(5279) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM1(5279))))  severity failure;
	assert RAM1(5280) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM1(5280))))  severity failure;
	assert RAM1(5281) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM1(5281))))  severity failure;
	assert RAM1(5282) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM1(5282))))  severity failure;
	assert RAM1(5283) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM1(5283))))  severity failure;
	assert RAM1(5284) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM1(5284))))  severity failure;
	assert RAM1(5285) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM1(5285))))  severity failure;
	assert RAM1(5286) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM1(5286))))  severity failure;
	assert RAM1(5287) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM1(5287))))  severity failure;
	assert RAM1(5288) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM1(5288))))  severity failure;
	assert RAM1(5289) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM1(5289))))  severity failure;
	assert RAM1(5290) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM1(5290))))  severity failure;
	assert RAM1(5291) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM1(5291))))  severity failure;
	assert RAM1(5292) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM1(5292))))  severity failure;
	assert RAM1(5293) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM1(5293))))  severity failure;
	assert RAM1(5294) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM1(5294))))  severity failure;
	assert RAM1(5295) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM1(5295))))  severity failure;
	assert RAM1(5296) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM1(5296))))  severity failure;
	assert RAM1(5297) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM1(5297))))  severity failure;
	assert RAM1(5298) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM1(5298))))  severity failure;
	assert RAM1(5299) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM1(5299))))  severity failure;
	assert RAM1(5300) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM1(5300))))  severity failure;
	assert RAM1(5301) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM1(5301))))  severity failure;
	assert RAM1(5302) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM1(5302))))  severity failure;
	assert RAM1(5303) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM1(5303))))  severity failure;
	assert RAM1(5304) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM1(5304))))  severity failure;
	assert RAM1(5305) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM1(5305))))  severity failure;
	assert RAM1(5306) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM1(5306))))  severity failure;
	assert RAM1(5307) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM1(5307))))  severity failure;
	assert RAM1(5308) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM1(5308))))  severity failure;
	assert RAM1(5309) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM1(5309))))  severity failure;
	assert RAM1(5310) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM1(5310))))  severity failure;
	assert RAM1(5311) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM1(5311))))  severity failure;
	assert RAM1(5312) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM1(5312))))  severity failure;
	assert RAM1(5313) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM1(5313))))  severity failure;
	assert RAM1(5314) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM1(5314))))  severity failure;
	assert RAM1(5315) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM1(5315))))  severity failure;
	assert RAM1(5316) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM1(5316))))  severity failure;
	assert RAM1(5317) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM1(5317))))  severity failure;
	assert RAM1(5318) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM1(5318))))  severity failure;
	assert RAM1(5319) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM1(5319))))  severity failure;
	assert RAM1(5320) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM1(5320))))  severity failure;
	assert RAM1(5321) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM1(5321))))  severity failure;
	assert RAM1(5322) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM1(5322))))  severity failure;
	assert RAM1(5323) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM1(5323))))  severity failure;
	assert RAM1(5324) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM1(5324))))  severity failure;
	assert RAM1(5325) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM1(5325))))  severity failure;
	assert RAM1(5326) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM1(5326))))  severity failure;
	assert RAM1(5327) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM1(5327))))  severity failure;
	assert RAM1(5328) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM1(5328))))  severity failure;
	assert RAM1(5329) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM1(5329))))  severity failure;
	assert RAM1(5330) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM1(5330))))  severity failure;
	assert RAM1(5331) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM1(5331))))  severity failure;
	assert RAM1(5332) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM1(5332))))  severity failure;
	assert RAM1(5333) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM1(5333))))  severity failure;
	assert RAM1(5334) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM1(5334))))  severity failure;
	assert RAM1(5335) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM1(5335))))  severity failure;
	assert RAM1(5336) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM1(5336))))  severity failure;
	assert RAM1(5337) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM1(5337))))  severity failure;
	assert RAM1(5338) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM1(5338))))  severity failure;
	assert RAM1(5339) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM1(5339))))  severity failure;
	assert RAM1(5340) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM1(5340))))  severity failure;
	assert RAM1(5341) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM1(5341))))  severity failure;
	assert RAM1(5342) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM1(5342))))  severity failure;
	assert RAM1(5343) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM1(5343))))  severity failure;
	assert RAM1(5344) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM1(5344))))  severity failure;
	assert RAM1(5345) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM1(5345))))  severity failure;
	assert RAM1(5346) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM1(5346))))  severity failure;
	assert RAM1(5347) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM1(5347))))  severity failure;
	assert RAM1(5348) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM1(5348))))  severity failure;
	assert RAM1(5349) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM1(5349))))  severity failure;
	assert RAM1(5350) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM1(5350))))  severity failure;
	assert RAM1(5351) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM1(5351))))  severity failure;
	assert RAM1(5352) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM1(5352))))  severity failure;
	assert RAM1(5353) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM1(5353))))  severity failure;
	assert RAM1(5354) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM1(5354))))  severity failure;
	assert RAM1(5355) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM1(5355))))  severity failure;
	assert RAM1(5356) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM1(5356))))  severity failure;
	assert RAM1(5357) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM1(5357))))  severity failure;
	assert RAM1(5358) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM1(5358))))  severity failure;
	assert RAM1(5359) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM1(5359))))  severity failure;
	assert RAM1(5360) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM1(5360))))  severity failure;
	assert RAM1(5361) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM1(5361))))  severity failure;
	assert RAM1(5362) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM1(5362))))  severity failure;
	assert RAM1(5363) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM1(5363))))  severity failure;
	assert RAM1(5364) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM1(5364))))  severity failure;
	assert RAM1(5365) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM1(5365))))  severity failure;
	assert RAM1(5366) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM1(5366))))  severity failure;
	assert RAM1(5367) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM1(5367))))  severity failure;
	assert RAM1(5368) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM1(5368))))  severity failure;
	assert RAM1(5369) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM1(5369))))  severity failure;
	assert RAM1(5370) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM1(5370))))  severity failure;
	assert RAM1(5371) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM1(5371))))  severity failure;
	assert RAM1(5372) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM1(5372))))  severity failure;
	assert RAM1(5373) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM1(5373))))  severity failure;
	assert RAM1(5374) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM1(5374))))  severity failure;
	assert RAM1(5375) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM1(5375))))  severity failure;
	assert RAM1(5376) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM1(5376))))  severity failure;
	assert RAM1(5377) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM1(5377))))  severity failure;
	assert RAM1(5378) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM1(5378))))  severity failure;
	assert RAM1(5379) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM1(5379))))  severity failure;
	assert RAM1(5380) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM1(5380))))  severity failure;
	assert RAM1(5381) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM1(5381))))  severity failure;
	assert RAM1(5382) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM1(5382))))  severity failure;
	assert RAM1(5383) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM1(5383))))  severity failure;
	assert RAM1(5384) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM1(5384))))  severity failure;
	assert RAM1(5385) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM1(5385))))  severity failure;
	assert RAM1(5386) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM1(5386))))  severity failure;
	assert RAM1(5387) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM1(5387))))  severity failure;
	assert RAM1(5388) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM1(5388))))  severity failure;
	assert RAM1(5389) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM1(5389))))  severity failure;
	assert RAM1(5390) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM1(5390))))  severity failure;
	assert RAM1(5391) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM1(5391))))  severity failure;
	assert RAM1(5392) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM1(5392))))  severity failure;
	assert RAM1(5393) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM1(5393))))  severity failure;
	assert RAM1(5394) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM1(5394))))  severity failure;
	assert RAM1(5395) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM1(5395))))  severity failure;
	assert RAM1(5396) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM1(5396))))  severity failure;
	assert RAM1(5397) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM1(5397))))  severity failure;
	assert RAM1(5398) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM1(5398))))  severity failure;
	assert RAM1(5399) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM1(5399))))  severity failure;
	assert RAM1(5400) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM1(5400))))  severity failure;
	assert RAM1(5401) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM1(5401))))  severity failure;
	assert RAM1(5402) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM1(5402))))  severity failure;
	assert RAM1(5403) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM1(5403))))  severity failure;
	assert RAM1(5404) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM1(5404))))  severity failure;
	assert RAM1(5405) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM1(5405))))  severity failure;
	assert RAM1(5406) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM1(5406))))  severity failure;
	assert RAM1(5407) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM1(5407))))  severity failure;
	assert RAM1(5408) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM1(5408))))  severity failure;
	assert RAM1(5409) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM1(5409))))  severity failure;
	assert RAM1(5410) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM1(5410))))  severity failure;
	assert RAM1(5411) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM1(5411))))  severity failure;
	assert RAM1(5412) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM1(5412))))  severity failure;
	assert RAM1(5413) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM1(5413))))  severity failure;
	assert RAM1(5414) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM1(5414))))  severity failure;
	assert RAM1(5415) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM1(5415))))  severity failure;
	assert RAM1(5416) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM1(5416))))  severity failure;
	assert RAM1(5417) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM1(5417))))  severity failure;
	assert RAM1(5418) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM1(5418))))  severity failure;
	assert RAM1(5419) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM1(5419))))  severity failure;
	assert RAM1(5420) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM1(5420))))  severity failure;
	assert RAM1(5421) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM1(5421))))  severity failure;
	assert RAM1(5422) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM1(5422))))  severity failure;
	assert RAM1(5423) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM1(5423))))  severity failure;
	assert RAM1(5424) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM1(5424))))  severity failure;
	assert RAM1(5425) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM1(5425))))  severity failure;
	assert RAM1(5426) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM1(5426))))  severity failure;
	assert RAM1(5427) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM1(5427))))  severity failure;
	assert RAM1(5428) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM1(5428))))  severity failure;
	assert RAM1(5429) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM1(5429))))  severity failure;
	assert RAM1(5430) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM1(5430))))  severity failure;
	assert RAM1(5431) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM1(5431))))  severity failure;
	assert RAM1(5432) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM1(5432))))  severity failure;
	assert RAM1(5433) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM1(5433))))  severity failure;
	assert RAM1(5434) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM1(5434))))  severity failure;
	assert RAM1(5435) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM1(5435))))  severity failure;
	assert RAM1(5436) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM1(5436))))  severity failure;
	assert RAM1(5437) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM1(5437))))  severity failure;
	assert RAM1(5438) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM1(5438))))  severity failure;
	assert RAM1(5439) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM1(5439))))  severity failure;
	assert RAM1(5440) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM1(5440))))  severity failure;
	assert RAM1(5441) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM1(5441))))  severity failure;
	assert RAM1(5442) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM1(5442))))  severity failure;
	assert RAM1(5443) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM1(5443))))  severity failure;
	assert RAM1(5444) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM1(5444))))  severity failure;
	assert RAM1(5445) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM1(5445))))  severity failure;
	assert RAM1(5446) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM1(5446))))  severity failure;
	assert RAM1(5447) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM1(5447))))  severity failure;
	assert RAM1(5448) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM1(5448))))  severity failure;
	assert RAM1(5449) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM1(5449))))  severity failure;
	assert RAM1(5450) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM1(5450))))  severity failure;
	assert RAM1(5451) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM1(5451))))  severity failure;
	assert RAM1(5452) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM1(5452))))  severity failure;
	assert RAM1(5453) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM1(5453))))  severity failure;
	assert RAM1(5454) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM1(5454))))  severity failure;
	assert RAM1(5455) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM1(5455))))  severity failure;
	assert RAM1(5456) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM1(5456))))  severity failure;
	assert RAM1(5457) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM1(5457))))  severity failure;
	assert RAM1(5458) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM1(5458))))  severity failure;
	assert RAM1(5459) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM1(5459))))  severity failure;
	assert RAM1(5460) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM1(5460))))  severity failure;
	assert RAM1(5461) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM1(5461))))  severity failure;
	assert RAM1(5462) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM1(5462))))  severity failure;
	assert RAM1(5463) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM1(5463))))  severity failure;
	assert RAM1(5464) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM1(5464))))  severity failure;
	assert RAM1(5465) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM1(5465))))  severity failure;
	assert RAM1(5466) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM1(5466))))  severity failure;
	assert RAM1(5467) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM1(5467))))  severity failure;
	assert RAM1(5468) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM1(5468))))  severity failure;
	assert RAM1(5469) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM1(5469))))  severity failure;
	assert RAM1(5470) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM1(5470))))  severity failure;
	assert RAM1(5471) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM1(5471))))  severity failure;
	assert RAM1(5472) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM1(5472))))  severity failure;
	assert RAM1(5473) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM1(5473))))  severity failure;
	assert RAM1(5474) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM1(5474))))  severity failure;
	assert RAM1(5475) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM1(5475))))  severity failure;
	assert RAM1(5476) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM1(5476))))  severity failure;
	assert RAM1(5477) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM1(5477))))  severity failure;
	assert RAM1(5478) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM1(5478))))  severity failure;
	assert RAM1(5479) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM1(5479))))  severity failure;
	assert RAM1(5480) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM1(5480))))  severity failure;
	assert RAM1(5481) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM1(5481))))  severity failure;
	assert RAM1(5482) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM1(5482))))  severity failure;
	assert RAM1(5483) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM1(5483))))  severity failure;
	assert RAM1(5484) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM1(5484))))  severity failure;
	assert RAM1(5485) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM1(5485))))  severity failure;
	assert RAM1(5486) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM1(5486))))  severity failure;
	assert RAM1(5487) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM1(5487))))  severity failure;
	assert RAM1(5488) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM1(5488))))  severity failure;
	assert RAM1(5489) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM1(5489))))  severity failure;
	assert RAM1(5490) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM1(5490))))  severity failure;
	assert RAM1(5491) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM1(5491))))  severity failure;
	assert RAM1(5492) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM1(5492))))  severity failure;
	assert RAM1(5493) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM1(5493))))  severity failure;
	assert RAM1(5494) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM1(5494))))  severity failure;
	assert RAM1(5495) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM1(5495))))  severity failure;
	assert RAM1(5496) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM1(5496))))  severity failure;
	assert RAM1(5497) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM1(5497))))  severity failure;
	assert RAM1(5498) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM1(5498))))  severity failure;
	assert RAM1(5499) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM1(5499))))  severity failure;
	assert RAM1(5500) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM1(5500))))  severity failure;
	assert RAM1(5501) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM1(5501))))  severity failure;
	assert RAM1(5502) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM1(5502))))  severity failure;
	assert RAM1(5503) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM1(5503))))  severity failure;
	assert RAM1(5504) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM1(5504))))  severity failure;
	assert RAM1(5505) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM1(5505))))  severity failure;
	assert RAM1(5506) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM1(5506))))  severity failure;
	assert RAM1(5507) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM1(5507))))  severity failure;
	assert RAM1(5508) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM1(5508))))  severity failure;
	assert RAM1(5509) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM1(5509))))  severity failure;
	assert RAM1(5510) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM1(5510))))  severity failure;
	assert RAM1(5511) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM1(5511))))  severity failure;
	assert RAM1(5512) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM1(5512))))  severity failure;
	assert RAM1(5513) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM1(5513))))  severity failure;
	assert RAM1(5514) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM1(5514))))  severity failure;
	assert RAM1(5515) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM1(5515))))  severity failure;
	assert RAM1(5516) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM1(5516))))  severity failure;
	assert RAM1(5517) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM1(5517))))  severity failure;
	assert RAM1(5518) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM1(5518))))  severity failure;
	assert RAM1(5519) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM1(5519))))  severity failure;
	assert RAM1(5520) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM1(5520))))  severity failure;
	assert RAM1(5521) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM1(5521))))  severity failure;
	assert RAM1(5522) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM1(5522))))  severity failure;
	assert RAM1(5523) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM1(5523))))  severity failure;
	assert RAM1(5524) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM1(5524))))  severity failure;
	assert RAM1(5525) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM1(5525))))  severity failure;
	assert RAM1(5526) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM1(5526))))  severity failure;
	assert RAM1(5527) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM1(5527))))  severity failure;
	assert RAM1(5528) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM1(5528))))  severity failure;
	assert RAM1(5529) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM1(5529))))  severity failure;
	assert RAM1(5530) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM1(5530))))  severity failure;
	assert RAM1(5531) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM1(5531))))  severity failure;
	assert RAM1(5532) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM1(5532))))  severity failure;
	assert RAM1(5533) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM1(5533))))  severity failure;
	assert RAM1(5534) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM1(5534))))  severity failure;
	assert RAM1(5535) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM1(5535))))  severity failure;
	assert RAM1(5536) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM1(5536))))  severity failure;
	assert RAM1(5537) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM1(5537))))  severity failure;
	assert RAM1(5538) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM1(5538))))  severity failure;
	assert RAM1(5539) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM1(5539))))  severity failure;
	assert RAM1(5540) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM1(5540))))  severity failure;
	assert RAM1(5541) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM1(5541))))  severity failure;
	assert RAM1(5542) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM1(5542))))  severity failure;
	assert RAM1(5543) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM1(5543))))  severity failure;
	assert RAM1(5544) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM1(5544))))  severity failure;
	assert RAM1(5545) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM1(5545))))  severity failure;
	assert RAM1(5546) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM1(5546))))  severity failure;
	assert RAM1(5547) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM1(5547))))  severity failure;
	assert RAM1(5548) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM1(5548))))  severity failure;
	assert RAM1(5549) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM1(5549))))  severity failure;
	assert RAM1(5550) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM1(5550))))  severity failure;
	assert RAM1(5551) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM1(5551))))  severity failure;
	assert RAM1(5552) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM1(5552))))  severity failure;
	assert RAM1(5553) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM1(5553))))  severity failure;
	assert RAM1(5554) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM1(5554))))  severity failure;
	assert RAM1(5555) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM1(5555))))  severity failure;
	assert RAM1(5556) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM1(5556))))  severity failure;
	assert RAM1(5557) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM1(5557))))  severity failure;
	assert RAM1(5558) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM1(5558))))  severity failure;
	assert RAM1(5559) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM1(5559))))  severity failure;
	assert RAM1(5560) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM1(5560))))  severity failure;
	assert RAM1(5561) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM1(5561))))  severity failure;
	assert RAM1(5562) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM1(5562))))  severity failure;
	assert RAM1(5563) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM1(5563))))  severity failure;
	assert RAM1(5564) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM1(5564))))  severity failure;
	assert RAM1(5565) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM1(5565))))  severity failure;
	assert RAM1(5566) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM1(5566))))  severity failure;
	assert RAM1(5567) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM1(5567))))  severity failure;
	assert RAM1(5568) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM1(5568))))  severity failure;
	assert RAM1(5569) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM1(5569))))  severity failure;
	assert RAM1(5570) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM1(5570))))  severity failure;
	assert RAM1(5571) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM1(5571))))  severity failure;
	assert RAM1(5572) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM1(5572))))  severity failure;
	assert RAM1(5573) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM1(5573))))  severity failure;
	assert RAM1(5574) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM1(5574))))  severity failure;
	assert RAM1(5575) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM1(5575))))  severity failure;
	assert RAM1(5576) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM1(5576))))  severity failure;
	assert RAM1(5577) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM1(5577))))  severity failure;
	assert RAM1(5578) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM1(5578))))  severity failure;
	assert RAM1(5579) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM1(5579))))  severity failure;
	assert RAM1(5580) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM1(5580))))  severity failure;
	assert RAM1(5581) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM1(5581))))  severity failure;
	assert RAM1(5582) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM1(5582))))  severity failure;
	assert RAM1(5583) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM1(5583))))  severity failure;
	assert RAM1(5584) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM1(5584))))  severity failure;
	assert RAM1(5585) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM1(5585))))  severity failure;
	assert RAM1(5586) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM1(5586))))  severity failure;
	assert RAM1(5587) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM1(5587))))  severity failure;
	assert RAM1(5588) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM1(5588))))  severity failure;
	assert RAM1(5589) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM1(5589))))  severity failure;
	assert RAM1(5590) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM1(5590))))  severity failure;
	assert RAM1(5591) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM1(5591))))  severity failure;
	assert RAM1(5592) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM1(5592))))  severity failure;
	assert RAM1(5593) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM1(5593))))  severity failure;
	assert RAM1(5594) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM1(5594))))  severity failure;
	assert RAM1(5595) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM1(5595))))  severity failure;
	assert RAM1(5596) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM1(5596))))  severity failure;
	assert RAM1(5597) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM1(5597))))  severity failure;
	assert RAM1(5598) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM1(5598))))  severity failure;
	assert RAM1(5599) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM1(5599))))  severity failure;
	assert RAM1(5600) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM1(5600))))  severity failure;
	assert RAM1(5601) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM1(5601))))  severity failure;
	assert RAM1(5602) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM1(5602))))  severity failure;
	assert RAM1(5603) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM1(5603))))  severity failure;
	assert RAM1(5604) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM1(5604))))  severity failure;
	assert RAM1(5605) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM1(5605))))  severity failure;
	assert RAM1(5606) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM1(5606))))  severity failure;
	assert RAM1(5607) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM1(5607))))  severity failure;
	assert RAM1(5608) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM1(5608))))  severity failure;
	assert RAM1(5609) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM1(5609))))  severity failure;
	assert RAM1(5610) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM1(5610))))  severity failure;
	assert RAM1(5611) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM1(5611))))  severity failure;
	assert RAM1(5612) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM1(5612))))  severity failure;
	assert RAM1(5613) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM1(5613))))  severity failure;
	assert RAM1(5614) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM1(5614))))  severity failure;
	assert RAM1(5615) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM1(5615))))  severity failure;
	assert RAM1(5616) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM1(5616))))  severity failure;
	assert RAM1(5617) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM1(5617))))  severity failure;
	assert RAM1(5618) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM1(5618))))  severity failure;
	assert RAM1(5619) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM1(5619))))  severity failure;
	assert RAM1(5620) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM1(5620))))  severity failure;
	assert RAM1(5621) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM1(5621))))  severity failure;
	assert RAM1(5622) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM1(5622))))  severity failure;
	assert RAM1(5623) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM1(5623))))  severity failure;
	assert RAM1(5624) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM1(5624))))  severity failure;
	assert RAM1(5625) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM1(5625))))  severity failure;
	assert RAM1(5626) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM1(5626))))  severity failure;
	assert RAM1(5627) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM1(5627))))  severity failure;
	assert RAM1(5628) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM1(5628))))  severity failure;
	assert RAM1(5629) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM1(5629))))  severity failure;
	assert RAM1(5630) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM1(5630))))  severity failure;
	assert RAM1(5631) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM1(5631))))  severity failure;
	assert RAM1(5632) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM1(5632))))  severity failure;
	assert RAM1(5633) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM1(5633))))  severity failure;
	assert RAM1(5634) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM1(5634))))  severity failure;
	assert RAM1(5635) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM1(5635))))  severity failure;
	assert RAM1(5636) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM1(5636))))  severity failure;
	assert RAM1(5637) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM1(5637))))  severity failure;
	assert RAM1(5638) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM1(5638))))  severity failure;
	assert RAM1(5639) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM1(5639))))  severity failure;
	assert RAM1(5640) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM1(5640))))  severity failure;
	assert RAM1(5641) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM1(5641))))  severity failure;
	assert RAM1(5642) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM1(5642))))  severity failure;
	assert RAM1(5643) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM1(5643))))  severity failure;
	assert RAM1(5644) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM1(5644))))  severity failure;
	assert RAM1(5645) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM1(5645))))  severity failure;
	assert RAM1(5646) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM1(5646))))  severity failure;
	assert RAM1(5647) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM1(5647))))  severity failure;
	assert RAM1(5648) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM1(5648))))  severity failure;
	assert RAM1(5649) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM1(5649))))  severity failure;
	assert RAM1(5650) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM1(5650))))  severity failure;
	assert RAM1(5651) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM1(5651))))  severity failure;
	assert RAM1(5652) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM1(5652))))  severity failure;
	assert RAM1(5653) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM1(5653))))  severity failure;
	assert RAM1(5654) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM1(5654))))  severity failure;
	assert RAM1(5655) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM1(5655))))  severity failure;
	assert RAM1(5656) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM1(5656))))  severity failure;
	assert RAM1(5657) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM1(5657))))  severity failure;
	assert RAM1(5658) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM1(5658))))  severity failure;
	assert RAM1(5659) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM1(5659))))  severity failure;
	assert RAM1(5660) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM1(5660))))  severity failure;
	assert RAM1(5661) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM1(5661))))  severity failure;
	assert RAM1(5662) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM1(5662))))  severity failure;
	assert RAM1(5663) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM1(5663))))  severity failure;
	assert RAM1(5664) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM1(5664))))  severity failure;
	assert RAM1(5665) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM1(5665))))  severity failure;
	assert RAM1(5666) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM1(5666))))  severity failure;
	assert RAM1(5667) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM1(5667))))  severity failure;
	assert RAM1(5668) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM1(5668))))  severity failure;
	assert RAM1(5669) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM1(5669))))  severity failure;
	assert RAM1(5670) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM1(5670))))  severity failure;
	assert RAM1(5671) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM1(5671))))  severity failure;
	assert RAM1(5672) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM1(5672))))  severity failure;
	assert RAM1(5673) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM1(5673))))  severity failure;
	assert RAM1(5674) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM1(5674))))  severity failure;
	assert RAM1(5675) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM1(5675))))  severity failure;
	assert RAM1(5676) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM1(5676))))  severity failure;
	assert RAM1(5677) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM1(5677))))  severity failure;
	assert RAM1(5678) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM1(5678))))  severity failure;
	assert RAM1(5679) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM1(5679))))  severity failure;
	assert RAM1(5680) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM1(5680))))  severity failure;
	assert RAM1(5681) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM1(5681))))  severity failure;
	assert RAM1(5682) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM1(5682))))  severity failure;
	assert RAM1(5683) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM1(5683))))  severity failure;
	assert RAM1(5684) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM1(5684))))  severity failure;
	assert RAM1(5685) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM1(5685))))  severity failure;
	assert RAM1(5686) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM1(5686))))  severity failure;
	assert RAM1(5687) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM1(5687))))  severity failure;
	assert RAM1(5688) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM1(5688))))  severity failure;
	assert RAM1(5689) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM1(5689))))  severity failure;
	assert RAM1(5690) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM1(5690))))  severity failure;
	assert RAM1(5691) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM1(5691))))  severity failure;
	assert RAM1(5692) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM1(5692))))  severity failure;
	assert RAM1(5693) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM1(5693))))  severity failure;
	assert RAM1(5694) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM1(5694))))  severity failure;
	assert RAM1(5695) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM1(5695))))  severity failure;
	assert RAM1(5696) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM1(5696))))  severity failure;
	assert RAM1(5697) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM1(5697))))  severity failure;
	assert RAM1(5698) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM1(5698))))  severity failure;
	assert RAM1(5699) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM1(5699))))  severity failure;
	assert RAM1(5700) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM1(5700))))  severity failure;
	assert RAM1(5701) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM1(5701))))  severity failure;
	assert RAM1(5702) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM1(5702))))  severity failure;
	assert RAM1(5703) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM1(5703))))  severity failure;
	assert RAM1(5704) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM1(5704))))  severity failure;
	assert RAM1(5705) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM1(5705))))  severity failure;
	assert RAM1(5706) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM1(5706))))  severity failure;
	assert RAM1(5707) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM1(5707))))  severity failure;
	assert RAM1(5708) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM1(5708))))  severity failure;
	assert RAM1(5709) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM1(5709))))  severity failure;
	assert RAM1(5710) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM1(5710))))  severity failure;
	assert RAM1(5711) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM1(5711))))  severity failure;
	assert RAM1(5712) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM1(5712))))  severity failure;
	assert RAM1(5713) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM1(5713))))  severity failure;
	assert RAM1(5714) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM1(5714))))  severity failure;
	assert RAM1(5715) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM1(5715))))  severity failure;
	assert RAM1(5716) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM1(5716))))  severity failure;
	assert RAM1(5717) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM1(5717))))  severity failure;
	assert RAM1(5718) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM1(5718))))  severity failure;
	assert RAM1(5719) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM1(5719))))  severity failure;
	assert RAM1(5720) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM1(5720))))  severity failure;
	assert RAM1(5721) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM1(5721))))  severity failure;
	assert RAM1(5722) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM1(5722))))  severity failure;
	assert RAM1(5723) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM1(5723))))  severity failure;
	assert RAM1(5724) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM1(5724))))  severity failure;
	assert RAM1(5725) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM1(5725))))  severity failure;
	assert RAM1(5726) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM1(5726))))  severity failure;
	assert RAM1(5727) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM1(5727))))  severity failure;
	assert RAM1(5728) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM1(5728))))  severity failure;
	assert RAM1(5729) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM1(5729))))  severity failure;
	assert RAM1(5730) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM1(5730))))  severity failure;
	assert RAM1(5731) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM1(5731))))  severity failure;
	assert RAM1(5732) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM1(5732))))  severity failure;
	assert RAM1(5733) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM1(5733))))  severity failure;
	assert RAM1(5734) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM1(5734))))  severity failure;
	assert RAM1(5735) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM1(5735))))  severity failure;
	assert RAM1(5736) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM1(5736))))  severity failure;
	assert RAM1(5737) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM1(5737))))  severity failure;
	assert RAM1(5738) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM1(5738))))  severity failure;
	assert RAM1(5739) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM1(5739))))  severity failure;
	assert RAM1(5740) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM1(5740))))  severity failure;
	assert RAM1(5741) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM1(5741))))  severity failure;
	assert RAM1(5742) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM1(5742))))  severity failure;
	assert RAM1(5743) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM1(5743))))  severity failure;
	assert RAM1(5744) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM1(5744))))  severity failure;
	assert RAM1(5745) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM1(5745))))  severity failure;
	assert RAM1(5746) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM1(5746))))  severity failure;
	assert RAM1(5747) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM1(5747))))  severity failure;
	assert RAM1(5748) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM1(5748))))  severity failure;
	assert RAM1(5749) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM1(5749))))  severity failure;
	assert RAM1(5750) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM1(5750))))  severity failure;
	assert RAM1(5751) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM1(5751))))  severity failure;
	assert RAM1(5752) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM1(5752))))  severity failure;
	assert RAM1(5753) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM1(5753))))  severity failure;
	assert RAM1(5754) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM1(5754))))  severity failure;
	assert RAM1(5755) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM1(5755))))  severity failure;
	assert RAM1(5756) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM1(5756))))  severity failure;
	assert RAM1(5757) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM1(5757))))  severity failure;
	assert RAM1(5758) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM1(5758))))  severity failure;
	assert RAM1(5759) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM1(5759))))  severity failure;
	assert RAM1(5760) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM1(5760))))  severity failure;
	assert RAM1(5761) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM1(5761))))  severity failure;
	assert RAM1(5762) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM1(5762))))  severity failure;
	assert RAM1(5763) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM1(5763))))  severity failure;
	assert RAM1(5764) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM1(5764))))  severity failure;
	assert RAM1(5765) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM1(5765))))  severity failure;
	assert RAM1(5766) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM1(5766))))  severity failure;
	assert RAM1(5767) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM1(5767))))  severity failure;
	assert RAM1(5768) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM1(5768))))  severity failure;
	assert RAM1(5769) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM1(5769))))  severity failure;
	assert RAM1(5770) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM1(5770))))  severity failure;
	assert RAM1(5771) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM1(5771))))  severity failure;
	assert RAM1(5772) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM1(5772))))  severity failure;
	assert RAM1(5773) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM1(5773))))  severity failure;
	assert RAM1(5774) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM1(5774))))  severity failure;
	assert RAM1(5775) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM1(5775))))  severity failure;
	assert RAM1(5776) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM1(5776))))  severity failure;
	assert RAM1(5777) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM1(5777))))  severity failure;
	assert RAM1(5778) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM1(5778))))  severity failure;
	assert RAM1(5779) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM1(5779))))  severity failure;
	assert RAM1(5780) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM1(5780))))  severity failure;
	assert RAM1(5781) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM1(5781))))  severity failure;
	assert RAM1(5782) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM1(5782))))  severity failure;
	assert RAM1(5783) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM1(5783))))  severity failure;
	assert RAM1(5784) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM1(5784))))  severity failure;
	assert RAM1(5785) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM1(5785))))  severity failure;
	assert RAM1(5786) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM1(5786))))  severity failure;
	assert RAM1(5787) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM1(5787))))  severity failure;
	assert RAM1(5788) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM1(5788))))  severity failure;
	assert RAM1(5789) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM1(5789))))  severity failure;
	assert RAM1(5790) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM1(5790))))  severity failure;
	assert RAM1(5791) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM1(5791))))  severity failure;
	assert RAM1(5792) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM1(5792))))  severity failure;
	assert RAM1(5793) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM1(5793))))  severity failure;
	assert RAM1(5794) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM1(5794))))  severity failure;
	assert RAM1(5795) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM1(5795))))  severity failure;
	assert RAM1(5796) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM1(5796))))  severity failure;
	assert RAM1(5797) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM1(5797))))  severity failure;
	assert RAM1(5798) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM1(5798))))  severity failure;
	assert RAM1(5799) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM1(5799))))  severity failure;
	assert RAM1(5800) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM1(5800))))  severity failure;
	assert RAM1(5801) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM1(5801))))  severity failure;
	assert RAM1(5802) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM1(5802))))  severity failure;
	assert RAM1(5803) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM1(5803))))  severity failure;
	assert RAM1(5804) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM1(5804))))  severity failure;
	assert RAM1(5805) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM1(5805))))  severity failure;
	assert RAM1(5806) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM1(5806))))  severity failure;
	assert RAM1(5807) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM1(5807))))  severity failure;
	assert RAM1(5808) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM1(5808))))  severity failure;
	assert RAM1(5809) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM1(5809))))  severity failure;
	assert RAM1(5810) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM1(5810))))  severity failure;
	assert RAM1(5811) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM1(5811))))  severity failure;
	assert RAM1(5812) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM1(5812))))  severity failure;
	assert RAM1(5813) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM1(5813))))  severity failure;
	assert RAM1(5814) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM1(5814))))  severity failure;
	assert RAM1(5815) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM1(5815))))  severity failure;
	assert RAM1(5816) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM1(5816))))  severity failure;
	assert RAM1(5817) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM1(5817))))  severity failure;
	assert RAM1(5818) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM1(5818))))  severity failure;
	assert RAM1(5819) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM1(5819))))  severity failure;
	assert RAM1(5820) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM1(5820))))  severity failure;
	assert RAM1(5821) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM1(5821))))  severity failure;
	assert RAM1(5822) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM1(5822))))  severity failure;
	assert RAM1(5823) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM1(5823))))  severity failure;
	assert RAM1(5824) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM1(5824))))  severity failure;
	assert RAM1(5825) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM1(5825))))  severity failure;
	assert RAM1(5826) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM1(5826))))  severity failure;
	assert RAM1(5827) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM1(5827))))  severity failure;
	assert RAM1(5828) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM1(5828))))  severity failure;
	assert RAM1(5829) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM1(5829))))  severity failure;
	assert RAM1(5830) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM1(5830))))  severity failure;
	assert RAM1(5831) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM1(5831))))  severity failure;
	assert RAM1(5832) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM1(5832))))  severity failure;
	assert RAM1(5833) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM1(5833))))  severity failure;
	assert RAM1(5834) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM1(5834))))  severity failure;
	assert RAM1(5835) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM1(5835))))  severity failure;
	assert RAM1(5836) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM1(5836))))  severity failure;
	assert RAM1(5837) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM1(5837))))  severity failure;
	assert RAM1(5838) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM1(5838))))  severity failure;
	assert RAM1(5839) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM1(5839))))  severity failure;
	assert RAM1(5840) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM1(5840))))  severity failure;
	assert RAM1(5841) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM1(5841))))  severity failure;
	assert RAM1(5842) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM1(5842))))  severity failure;
	assert RAM1(5843) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM1(5843))))  severity failure;
	assert RAM1(5844) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM1(5844))))  severity failure;
	assert RAM1(5845) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM1(5845))))  severity failure;
	assert RAM1(5846) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM1(5846))))  severity failure;
	assert RAM1(5847) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM1(5847))))  severity failure;
	assert RAM1(5848) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM1(5848))))  severity failure;
	assert RAM1(5849) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM1(5849))))  severity failure;
	assert RAM1(5850) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM1(5850))))  severity failure;
	assert RAM1(5851) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM1(5851))))  severity failure;
	assert RAM1(5852) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM1(5852))))  severity failure;
	assert RAM1(5853) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM1(5853))))  severity failure;
	assert RAM1(5854) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM1(5854))))  severity failure;
	assert RAM1(5855) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM1(5855))))  severity failure;
	assert RAM1(5856) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM1(5856))))  severity failure;
	assert RAM1(5857) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM1(5857))))  severity failure;
	assert RAM1(5858) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM1(5858))))  severity failure;
	assert RAM1(5859) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM1(5859))))  severity failure;
	assert RAM1(5860) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM1(5860))))  severity failure;
	assert RAM1(5861) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM1(5861))))  severity failure;
	assert RAM1(5862) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM1(5862))))  severity failure;
	assert RAM1(5863) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM1(5863))))  severity failure;
	assert RAM1(5864) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM1(5864))))  severity failure;
	assert RAM1(5865) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM1(5865))))  severity failure;
	assert RAM1(5866) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM1(5866))))  severity failure;
	assert RAM1(5867) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM1(5867))))  severity failure;
	assert RAM1(5868) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM1(5868))))  severity failure;
	assert RAM1(5869) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM1(5869))))  severity failure;
	assert RAM1(5870) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM1(5870))))  severity failure;
	assert RAM1(5871) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM1(5871))))  severity failure;
	assert RAM1(5872) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM1(5872))))  severity failure;
	assert RAM1(5873) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM1(5873))))  severity failure;
	assert RAM1(5874) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM1(5874))))  severity failure;
	assert RAM1(5875) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM1(5875))))  severity failure;
	assert RAM1(5876) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM1(5876))))  severity failure;
	assert RAM1(5877) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM1(5877))))  severity failure;
	assert RAM1(5878) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM1(5878))))  severity failure;
	assert RAM1(5879) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM1(5879))))  severity failure;
	assert RAM1(5880) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM1(5880))))  severity failure;
	assert RAM1(5881) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM1(5881))))  severity failure;
	assert RAM1(5882) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM1(5882))))  severity failure;
	assert RAM1(5883) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM1(5883))))  severity failure;
	assert RAM1(5884) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM1(5884))))  severity failure;
	assert RAM1(5885) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM1(5885))))  severity failure;
	assert RAM1(5886) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM1(5886))))  severity failure;
	assert RAM1(5887) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM1(5887))))  severity failure;
	assert RAM1(5888) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM1(5888))))  severity failure;
	assert RAM1(5889) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM1(5889))))  severity failure;
	assert RAM1(5890) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM1(5890))))  severity failure;
	assert RAM1(5891) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM1(5891))))  severity failure;
	assert RAM1(5892) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM1(5892))))  severity failure;
	assert RAM1(5893) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM1(5893))))  severity failure;
	assert RAM1(5894) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM1(5894))))  severity failure;
	assert RAM1(5895) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM1(5895))))  severity failure;
	assert RAM1(5896) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM1(5896))))  severity failure;
	assert RAM1(5897) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM1(5897))))  severity failure;
	assert RAM1(5898) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM1(5898))))  severity failure;
	assert RAM1(5899) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM1(5899))))  severity failure;
	assert RAM1(5900) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM1(5900))))  severity failure;
	assert RAM1(5901) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM1(5901))))  severity failure;
	assert RAM1(5902) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM1(5902))))  severity failure;
	assert RAM1(5903) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM1(5903))))  severity failure;
	assert RAM1(5904) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM1(5904))))  severity failure;
	assert RAM1(5905) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM1(5905))))  severity failure;
	assert RAM1(5906) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM1(5906))))  severity failure;
	assert RAM1(5907) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM1(5907))))  severity failure;
	assert RAM1(5908) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM1(5908))))  severity failure;
	assert RAM1(5909) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM1(5909))))  severity failure;
	assert RAM1(5910) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM1(5910))))  severity failure;
	assert RAM1(5911) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM1(5911))))  severity failure;
	assert RAM1(5912) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM1(5912))))  severity failure;
	assert RAM1(5913) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM1(5913))))  severity failure;
	assert RAM1(5914) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM1(5914))))  severity failure;
	assert RAM1(5915) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM1(5915))))  severity failure;
	assert RAM1(5916) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM1(5916))))  severity failure;
	assert RAM1(5917) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM1(5917))))  severity failure;
	assert RAM1(5918) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM1(5918))))  severity failure;
	assert RAM1(5919) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM1(5919))))  severity failure;
	assert RAM1(5920) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM1(5920))))  severity failure;
	assert RAM1(5921) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM1(5921))))  severity failure;
	assert RAM1(5922) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM1(5922))))  severity failure;
	assert RAM1(5923) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM1(5923))))  severity failure;
	assert RAM1(5924) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM1(5924))))  severity failure;
	assert RAM1(5925) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM1(5925))))  severity failure;
	assert RAM1(5926) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM1(5926))))  severity failure;
	assert RAM1(5927) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM1(5927))))  severity failure;
	assert RAM1(5928) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM1(5928))))  severity failure;
	assert RAM1(5929) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM1(5929))))  severity failure;
	assert RAM1(5930) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM1(5930))))  severity failure;
	assert RAM1(5931) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM1(5931))))  severity failure;
	assert RAM1(5932) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM1(5932))))  severity failure;
	assert RAM1(5933) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM1(5933))))  severity failure;
	assert RAM1(5934) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM1(5934))))  severity failure;
	assert RAM1(5935) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM1(5935))))  severity failure;
	assert RAM1(5936) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM1(5936))))  severity failure;
	assert RAM1(5937) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM1(5937))))  severity failure;
	assert RAM1(5938) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM1(5938))))  severity failure;
	assert RAM1(5939) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM1(5939))))  severity failure;
	assert RAM1(5940) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM1(5940))))  severity failure;
	assert RAM1(5941) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM1(5941))))  severity failure;
	assert RAM1(5942) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM1(5942))))  severity failure;
	assert RAM1(5943) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM1(5943))))  severity failure;
	assert RAM1(5944) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM1(5944))))  severity failure;
	assert RAM1(5945) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM1(5945))))  severity failure;
	assert RAM1(5946) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM1(5946))))  severity failure;
	assert RAM1(5947) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM1(5947))))  severity failure;
	assert RAM1(5948) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM1(5948))))  severity failure;
	assert RAM1(5949) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM1(5949))))  severity failure;
	assert RAM1(5950) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM1(5950))))  severity failure;
	assert RAM1(5951) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM1(5951))))  severity failure;
	assert RAM1(5952) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM1(5952))))  severity failure;
	assert RAM1(5953) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM1(5953))))  severity failure;
	assert RAM1(5954) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM1(5954))))  severity failure;
	assert RAM1(5955) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM1(5955))))  severity failure;
	assert RAM1(5956) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM1(5956))))  severity failure;
	assert RAM1(5957) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM1(5957))))  severity failure;
	assert RAM1(5958) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM1(5958))))  severity failure;
	assert RAM1(5959) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM1(5959))))  severity failure;
	assert RAM1(5960) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM1(5960))))  severity failure;
	assert RAM1(5961) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM1(5961))))  severity failure;
	assert RAM1(5962) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM1(5962))))  severity failure;
	assert RAM1(5963) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM1(5963))))  severity failure;
	assert RAM1(5964) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM1(5964))))  severity failure;
	assert RAM1(5965) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM1(5965))))  severity failure;
	assert RAM1(5966) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM1(5966))))  severity failure;
	assert RAM1(5967) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM1(5967))))  severity failure;
	assert RAM1(5968) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM1(5968))))  severity failure;
	assert RAM1(5969) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM1(5969))))  severity failure;
	assert RAM1(5970) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM1(5970))))  severity failure;
	assert RAM1(5971) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM1(5971))))  severity failure;
	assert RAM1(5972) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM1(5972))))  severity failure;
	assert RAM1(5973) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM1(5973))))  severity failure;
	assert RAM1(5974) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM1(5974))))  severity failure;
	assert RAM1(5975) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM1(5975))))  severity failure;
	assert RAM1(5976) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM1(5976))))  severity failure;
	assert RAM1(5977) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM1(5977))))  severity failure;
	assert RAM1(5978) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM1(5978))))  severity failure;
	assert RAM1(5979) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM1(5979))))  severity failure;
	assert RAM1(5980) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM1(5980))))  severity failure;
	assert RAM1(5981) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM1(5981))))  severity failure;
	assert RAM1(5982) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM1(5982))))  severity failure;
	assert RAM1(5983) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM1(5983))))  severity failure;
	assert RAM1(5984) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM1(5984))))  severity failure;
	assert RAM1(5985) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM1(5985))))  severity failure;
	assert RAM1(5986) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM1(5986))))  severity failure;
	assert RAM1(5987) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM1(5987))))  severity failure;
	assert RAM1(5988) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM1(5988))))  severity failure;
	assert RAM1(5989) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM1(5989))))  severity failure;
	assert RAM1(5990) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM1(5990))))  severity failure;
	assert RAM1(5991) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM1(5991))))  severity failure;
	assert RAM1(5992) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM1(5992))))  severity failure;
	assert RAM1(5993) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM1(5993))))  severity failure;
	assert RAM1(5994) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM1(5994))))  severity failure;
	assert RAM1(5995) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM1(5995))))  severity failure;
	assert RAM1(5996) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM1(5996))))  severity failure;
	assert RAM1(5997) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM1(5997))))  severity failure;
	assert RAM1(5998) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM1(5998))))  severity failure;
	assert RAM1(5999) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM1(5999))))  severity failure;
	assert RAM1(6000) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM1(6000))))  severity failure;
	assert RAM1(6001) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM1(6001))))  severity failure;
	assert RAM1(6002) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM1(6002))))  severity failure;
	assert RAM1(6003) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM1(6003))))  severity failure;
	assert RAM1(6004) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM1(6004))))  severity failure;
	assert RAM1(6005) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM1(6005))))  severity failure;
	assert RAM1(6006) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM1(6006))))  severity failure;
	assert RAM1(6007) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM1(6007))))  severity failure;
	assert RAM1(6008) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM1(6008))))  severity failure;
	assert RAM1(6009) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM1(6009))))  severity failure;
	assert RAM1(6010) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM1(6010))))  severity failure;
	assert RAM1(6011) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM1(6011))))  severity failure;
	assert RAM1(6012) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM1(6012))))  severity failure;
	assert RAM1(6013) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM1(6013))))  severity failure;
	assert RAM1(6014) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM1(6014))))  severity failure;
	assert RAM1(6015) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM1(6015))))  severity failure;
	assert RAM1(6016) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM1(6016))))  severity failure;
	assert RAM1(6017) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM1(6017))))  severity failure;
	assert RAM1(6018) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM1(6018))))  severity failure;
	assert RAM1(6019) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM1(6019))))  severity failure;
	assert RAM1(6020) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM1(6020))))  severity failure;
	assert RAM1(6021) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM1(6021))))  severity failure;
	assert RAM1(6022) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM1(6022))))  severity failure;
	assert RAM1(6023) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM1(6023))))  severity failure;
	assert RAM1(6024) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM1(6024))))  severity failure;
	assert RAM1(6025) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM1(6025))))  severity failure;
	assert RAM1(6026) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM1(6026))))  severity failure;
	assert RAM1(6027) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM1(6027))))  severity failure;
	assert RAM1(6028) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM1(6028))))  severity failure;
	assert RAM1(6029) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM1(6029))))  severity failure;
	assert RAM1(6030) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM1(6030))))  severity failure;
	assert RAM1(6031) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM1(6031))))  severity failure;
	assert RAM1(6032) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM1(6032))))  severity failure;
	assert RAM1(6033) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM1(6033))))  severity failure;
	assert RAM1(6034) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM1(6034))))  severity failure;
	assert RAM1(6035) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM1(6035))))  severity failure;
	assert RAM1(6036) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM1(6036))))  severity failure;
	assert RAM1(6037) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM1(6037))))  severity failure;
	assert RAM1(6038) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM1(6038))))  severity failure;
	assert RAM1(6039) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM1(6039))))  severity failure;
	assert RAM1(6040) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM1(6040))))  severity failure;
	assert RAM1(6041) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM1(6041))))  severity failure;
	assert RAM1(6042) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM1(6042))))  severity failure;
	assert RAM1(6043) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM1(6043))))  severity failure;
	assert RAM1(6044) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM1(6044))))  severity failure;
	assert RAM1(6045) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM1(6045))))  severity failure;
	assert RAM1(6046) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM1(6046))))  severity failure;
	assert RAM1(6047) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM1(6047))))  severity failure;
	assert RAM1(6048) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM1(6048))))  severity failure;
	assert RAM1(6049) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM1(6049))))  severity failure;
	assert RAM1(6050) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM1(6050))))  severity failure;
	assert RAM1(6051) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM1(6051))))  severity failure;
	assert RAM1(6052) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM1(6052))))  severity failure;
	assert RAM1(6053) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM1(6053))))  severity failure;
	assert RAM1(6054) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM1(6054))))  severity failure;
	assert RAM1(6055) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM1(6055))))  severity failure;
	assert RAM1(6056) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM1(6056))))  severity failure;
	assert RAM1(6057) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM1(6057))))  severity failure;
	assert RAM1(6058) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM1(6058))))  severity failure;
	assert RAM1(6059) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM1(6059))))  severity failure;
	assert RAM1(6060) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM1(6060))))  severity failure;
	assert RAM1(6061) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM1(6061))))  severity failure;
	assert RAM1(6062) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM1(6062))))  severity failure;
	assert RAM1(6063) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM1(6063))))  severity failure;
	assert RAM1(6064) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM1(6064))))  severity failure;
	assert RAM1(6065) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM1(6065))))  severity failure;
	assert RAM1(6066) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM1(6066))))  severity failure;
	assert RAM1(6067) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM1(6067))))  severity failure;
	assert RAM1(6068) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM1(6068))))  severity failure;
	assert RAM1(6069) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM1(6069))))  severity failure;
	assert RAM1(6070) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM1(6070))))  severity failure;
	assert RAM1(6071) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM1(6071))))  severity failure;
	assert RAM1(6072) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM1(6072))))  severity failure;
	assert RAM1(6073) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM1(6073))))  severity failure;
	assert RAM1(6074) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM1(6074))))  severity failure;
	assert RAM1(6075) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM1(6075))))  severity failure;
	assert RAM1(6076) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM1(6076))))  severity failure;
	assert RAM1(6077) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM1(6077))))  severity failure;
	assert RAM1(6078) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM1(6078))))  severity failure;
	assert RAM1(6079) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM1(6079))))  severity failure;
	assert RAM1(6080) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM1(6080))))  severity failure;
	assert RAM1(6081) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM1(6081))))  severity failure;
	assert RAM1(6082) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM1(6082))))  severity failure;
	assert RAM1(6083) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM1(6083))))  severity failure;
	assert RAM1(6084) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM1(6084))))  severity failure;
	assert RAM1(6085) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM1(6085))))  severity failure;
	assert RAM1(6086) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM1(6086))))  severity failure;
	assert RAM1(6087) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM1(6087))))  severity failure;
	assert RAM1(6088) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM1(6088))))  severity failure;
	assert RAM1(6089) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM1(6089))))  severity failure;
	assert RAM1(6090) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM1(6090))))  severity failure;
	assert RAM1(6091) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM1(6091))))  severity failure;
	assert RAM1(6092) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM1(6092))))  severity failure;
	assert RAM1(6093) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM1(6093))))  severity failure;
	assert RAM1(6094) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM1(6094))))  severity failure;
	assert RAM1(6095) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM1(6095))))  severity failure;
	assert RAM1(6096) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM1(6096))))  severity failure;
	assert RAM1(6097) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM1(6097))))  severity failure;
	assert RAM1(6098) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM1(6098))))  severity failure;
	assert RAM1(6099) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM1(6099))))  severity failure;
	assert RAM1(6100) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM1(6100))))  severity failure;
	assert RAM1(6101) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM1(6101))))  severity failure;
	assert RAM1(6102) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM1(6102))))  severity failure;
	assert RAM1(6103) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM1(6103))))  severity failure;
	assert RAM1(6104) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM1(6104))))  severity failure;
	assert RAM1(6105) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM1(6105))))  severity failure;
	assert RAM1(6106) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM1(6106))))  severity failure;
	assert RAM1(6107) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM1(6107))))  severity failure;
	assert RAM1(6108) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM1(6108))))  severity failure;
	assert RAM1(6109) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM1(6109))))  severity failure;
	assert RAM1(6110) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM1(6110))))  severity failure;
	assert RAM1(6111) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM1(6111))))  severity failure;
	assert RAM1(6112) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM1(6112))))  severity failure;
	assert RAM1(6113) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM1(6113))))  severity failure;
	assert RAM1(6114) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM1(6114))))  severity failure;
	assert RAM1(6115) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM1(6115))))  severity failure;
	assert RAM1(6116) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM1(6116))))  severity failure;
	assert RAM1(6117) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM1(6117))))  severity failure;
	assert RAM1(6118) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM1(6118))))  severity failure;
	assert RAM1(6119) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM1(6119))))  severity failure;
	assert RAM1(6120) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM1(6120))))  severity failure;
	assert RAM1(6121) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM1(6121))))  severity failure;
	assert RAM1(6122) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM1(6122))))  severity failure;
	assert RAM1(6123) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM1(6123))))  severity failure;
	assert RAM1(6124) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM1(6124))))  severity failure;
	assert RAM1(6125) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM1(6125))))  severity failure;
	assert RAM1(6126) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM1(6126))))  severity failure;
	assert RAM1(6127) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM1(6127))))  severity failure;
	assert RAM1(6128) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM1(6128))))  severity failure;
	assert RAM1(6129) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM1(6129))))  severity failure;
	assert RAM1(6130) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM1(6130))))  severity failure;
	assert RAM1(6131) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM1(6131))))  severity failure;
	assert RAM1(6132) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM1(6132))))  severity failure;
	assert RAM1(6133) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM1(6133))))  severity failure;
	assert RAM1(6134) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM1(6134))))  severity failure;
	assert RAM1(6135) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM1(6135))))  severity failure;
	assert RAM1(6136) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM1(6136))))  severity failure;
	assert RAM1(6137) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM1(6137))))  severity failure;
	assert RAM1(6138) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM1(6138))))  severity failure;
	assert RAM1(6139) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM1(6139))))  severity failure;
	assert RAM1(6140) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM1(6140))))  severity failure;
	assert RAM1(6141) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM1(6141))))  severity failure;
	assert RAM1(6142) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM1(6142))))  severity failure;
	assert RAM1(6143) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM1(6143))))  severity failure;
	assert RAM1(6144) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM1(6144))))  severity failure;
	assert RAM1(6145) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM1(6145))))  severity failure;
	assert RAM1(6146) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM1(6146))))  severity failure;
	assert RAM1(6147) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM1(6147))))  severity failure;
	assert RAM1(6148) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM1(6148))))  severity failure;
	assert RAM1(6149) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM1(6149))))  severity failure;
	assert RAM1(6150) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM1(6150))))  severity failure;
	assert RAM1(6151) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM1(6151))))  severity failure;
	assert RAM1(6152) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM1(6152))))  severity failure;
	assert RAM1(6153) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM1(6153))))  severity failure;
	assert RAM1(6154) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM1(6154))))  severity failure;
	assert RAM1(6155) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM1(6155))))  severity failure;
	assert RAM1(6156) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM1(6156))))  severity failure;
	assert RAM1(6157) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM1(6157))))  severity failure;
	assert RAM1(6158) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM1(6158))))  severity failure;
	assert RAM1(6159) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM1(6159))))  severity failure;
	assert RAM1(6160) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM1(6160))))  severity failure;
	assert RAM1(6161) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM1(6161))))  severity failure;
	assert RAM1(6162) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM1(6162))))  severity failure;
	assert RAM1(6163) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM1(6163))))  severity failure;
	assert RAM1(6164) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM1(6164))))  severity failure;
	assert RAM1(6165) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM1(6165))))  severity failure;
	assert RAM1(6166) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM1(6166))))  severity failure;
	assert RAM1(6167) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM1(6167))))  severity failure;
	assert RAM1(6168) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM1(6168))))  severity failure;
	assert RAM1(6169) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM1(6169))))  severity failure;
	assert RAM1(6170) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM1(6170))))  severity failure;
	assert RAM1(6171) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM1(6171))))  severity failure;
	assert RAM1(6172) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM1(6172))))  severity failure;
	assert RAM1(6173) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM1(6173))))  severity failure;
	assert RAM1(6174) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM1(6174))))  severity failure;
	assert RAM1(6175) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM1(6175))))  severity failure;
	assert RAM1(6176) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM1(6176))))  severity failure;
	assert RAM1(6177) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM1(6177))))  severity failure;
	assert RAM1(6178) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM1(6178))))  severity failure;
	assert RAM1(6179) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM1(6179))))  severity failure;
	assert RAM1(6180) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM1(6180))))  severity failure;
	assert RAM1(6181) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM1(6181))))  severity failure;
	assert RAM1(6182) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM1(6182))))  severity failure;
	assert RAM1(6183) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM1(6183))))  severity failure;
	assert RAM1(6184) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM1(6184))))  severity failure;
	assert RAM1(6185) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM1(6185))))  severity failure;
	assert RAM1(6186) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM1(6186))))  severity failure;
	assert RAM1(6187) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM1(6187))))  severity failure;
	assert RAM1(6188) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM1(6188))))  severity failure;
	assert RAM1(6189) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM1(6189))))  severity failure;
	assert RAM1(6190) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM1(6190))))  severity failure;
	assert RAM1(6191) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM1(6191))))  severity failure;
	assert RAM1(6192) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM1(6192))))  severity failure;
	assert RAM1(6193) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM1(6193))))  severity failure;
	assert RAM1(6194) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM1(6194))))  severity failure;
	assert RAM1(6195) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM1(6195))))  severity failure;
	assert RAM1(6196) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM1(6196))))  severity failure;
	assert RAM1(6197) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM1(6197))))  severity failure;
	assert RAM1(6198) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM1(6198))))  severity failure;
	assert RAM1(6199) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM1(6199))))  severity failure;
	assert RAM1(6200) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM1(6200))))  severity failure;
	assert RAM1(6201) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM1(6201))))  severity failure;
	assert RAM1(6202) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM1(6202))))  severity failure;
	assert RAM1(6203) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM1(6203))))  severity failure;
	assert RAM1(6204) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM1(6204))))  severity failure;
	assert RAM1(6205) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM1(6205))))  severity failure;
	assert RAM1(6206) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM1(6206))))  severity failure;
	assert RAM1(6207) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM1(6207))))  severity failure;
	assert RAM1(6208) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM1(6208))))  severity failure;
	assert RAM1(6209) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM1(6209))))  severity failure;
	assert RAM1(6210) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM1(6210))))  severity failure;
	assert RAM1(6211) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM1(6211))))  severity failure;
	assert RAM1(6212) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM1(6212))))  severity failure;
	assert RAM1(6213) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM1(6213))))  severity failure;
	assert RAM1(6214) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM1(6214))))  severity failure;
	assert RAM1(6215) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM1(6215))))  severity failure;
	assert RAM1(6216) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM1(6216))))  severity failure;
	assert RAM1(6217) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM1(6217))))  severity failure;
	assert RAM1(6218) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM1(6218))))  severity failure;
	assert RAM1(6219) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM1(6219))))  severity failure;
	assert RAM1(6220) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM1(6220))))  severity failure;
	assert RAM1(6221) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM1(6221))))  severity failure;
	assert RAM1(6222) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM1(6222))))  severity failure;
	assert RAM1(6223) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM1(6223))))  severity failure;
	assert RAM1(6224) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM1(6224))))  severity failure;
	assert RAM1(6225) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM1(6225))))  severity failure;
	assert RAM1(6226) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM1(6226))))  severity failure;
	assert RAM1(6227) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM1(6227))))  severity failure;
	assert RAM1(6228) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM1(6228))))  severity failure;
	assert RAM1(6229) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM1(6229))))  severity failure;
	assert RAM1(6230) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM1(6230))))  severity failure;
	assert RAM1(6231) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM1(6231))))  severity failure;
	assert RAM1(6232) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM1(6232))))  severity failure;
	assert RAM1(6233) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM1(6233))))  severity failure;
	assert RAM1(6234) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM1(6234))))  severity failure;
	assert RAM1(6235) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM1(6235))))  severity failure;
	assert RAM1(6236) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM1(6236))))  severity failure;
	assert RAM1(6237) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM1(6237))))  severity failure;
	assert RAM1(6238) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM1(6238))))  severity failure;
	assert RAM1(6239) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM1(6239))))  severity failure;
	assert RAM1(6240) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM1(6240))))  severity failure;
	assert RAM1(6241) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM1(6241))))  severity failure;
	assert RAM1(6242) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM1(6242))))  severity failure;
	assert RAM1(6243) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM1(6243))))  severity failure;
	assert RAM1(6244) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM1(6244))))  severity failure;
	assert RAM1(6245) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM1(6245))))  severity failure;
	assert RAM1(6246) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM1(6246))))  severity failure;
	assert RAM1(6247) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM1(6247))))  severity failure;
	assert RAM1(6248) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM1(6248))))  severity failure;
	assert RAM1(6249) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM1(6249))))  severity failure;
	assert RAM1(6250) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM1(6250))))  severity failure;
	assert RAM1(6251) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM1(6251))))  severity failure;
	assert RAM1(6252) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM1(6252))))  severity failure;
	assert RAM1(6253) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM1(6253))))  severity failure;
	assert RAM1(6254) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM1(6254))))  severity failure;
	assert RAM1(6255) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM1(6255))))  severity failure;
	assert RAM1(6256) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM1(6256))))  severity failure;
	assert RAM1(6257) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM1(6257))))  severity failure;
	assert RAM1(6258) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM1(6258))))  severity failure;
	assert RAM1(6259) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM1(6259))))  severity failure;
	assert RAM1(6260) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM1(6260))))  severity failure;
	assert RAM1(6261) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM1(6261))))  severity failure;
	assert RAM1(6262) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM1(6262))))  severity failure;
	assert RAM1(6263) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM1(6263))))  severity failure;
	assert RAM1(6264) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM1(6264))))  severity failure;
	assert RAM1(6265) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM1(6265))))  severity failure;
	assert RAM1(6266) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM1(6266))))  severity failure;
	assert RAM1(6267) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM1(6267))))  severity failure;
	assert RAM1(6268) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM1(6268))))  severity failure;
	assert RAM1(6269) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM1(6269))))  severity failure;
	assert RAM1(6270) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM1(6270))))  severity failure;
	assert RAM1(6271) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM1(6271))))  severity failure;
	assert RAM1(6272) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM1(6272))))  severity failure;
	assert RAM1(6273) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM1(6273))))  severity failure;
	assert RAM1(6274) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM1(6274))))  severity failure;
	assert RAM1(6275) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM1(6275))))  severity failure;
	assert RAM1(6276) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM1(6276))))  severity failure;
	assert RAM1(6277) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM1(6277))))  severity failure;
	assert RAM1(6278) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM1(6278))))  severity failure;
	assert RAM1(6279) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM1(6279))))  severity failure;
	assert RAM1(6280) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM1(6280))))  severity failure;
	assert RAM1(6281) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM1(6281))))  severity failure;
	assert RAM1(6282) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM1(6282))))  severity failure;
	assert RAM1(6283) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM1(6283))))  severity failure;
	assert RAM1(6284) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM1(6284))))  severity failure;
	assert RAM1(6285) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM1(6285))))  severity failure;
	assert RAM1(6286) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM1(6286))))  severity failure;
	assert RAM1(6287) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM1(6287))))  severity failure;
	assert RAM1(6288) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM1(6288))))  severity failure;
	assert RAM1(6289) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM1(6289))))  severity failure;
	assert RAM1(6290) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM1(6290))))  severity failure;
	assert RAM1(6291) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM1(6291))))  severity failure;
	assert RAM1(6292) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM1(6292))))  severity failure;
	assert RAM1(6293) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM1(6293))))  severity failure;
	assert RAM1(6294) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM1(6294))))  severity failure;
	assert RAM1(6295) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM1(6295))))  severity failure;
	assert RAM1(6296) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM1(6296))))  severity failure;
	assert RAM1(6297) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM1(6297))))  severity failure;
	assert RAM1(6298) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM1(6298))))  severity failure;
	assert RAM1(6299) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM1(6299))))  severity failure;
	assert RAM1(6300) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM1(6300))))  severity failure;
	assert RAM1(6301) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM1(6301))))  severity failure;
	assert RAM1(6302) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM1(6302))))  severity failure;
	assert RAM1(6303) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM1(6303))))  severity failure;
	assert RAM1(6304) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM1(6304))))  severity failure;
	assert RAM1(6305) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM1(6305))))  severity failure;
	assert RAM1(6306) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM1(6306))))  severity failure;
	assert RAM1(6307) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM1(6307))))  severity failure;
	assert RAM1(6308) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM1(6308))))  severity failure;
	assert RAM1(6309) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM1(6309))))  severity failure;
	assert RAM1(6310) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM1(6310))))  severity failure;
	assert RAM1(6311) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM1(6311))))  severity failure;
	assert RAM1(6312) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM1(6312))))  severity failure;
	assert RAM1(6313) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM1(6313))))  severity failure;
	assert RAM1(6314) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM1(6314))))  severity failure;
	assert RAM1(6315) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM1(6315))))  severity failure;
	assert RAM1(6316) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM1(6316))))  severity failure;
	assert RAM1(6317) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM1(6317))))  severity failure;
	assert RAM1(6318) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM1(6318))))  severity failure;
	assert RAM1(6319) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM1(6319))))  severity failure;
	assert RAM1(6320) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM1(6320))))  severity failure;
	assert RAM1(6321) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM1(6321))))  severity failure;
	assert RAM1(6322) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM1(6322))))  severity failure;
	assert RAM1(6323) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM1(6323))))  severity failure;
	assert RAM1(6324) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM1(6324))))  severity failure;
	assert RAM1(6325) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM1(6325))))  severity failure;
	assert RAM1(6326) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM1(6326))))  severity failure;
	assert RAM1(6327) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM1(6327))))  severity failure;
	assert RAM1(6328) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM1(6328))))  severity failure;
	assert RAM1(6329) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM1(6329))))  severity failure;
	assert RAM1(6330) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM1(6330))))  severity failure;
	assert RAM1(6331) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM1(6331))))  severity failure;
	assert RAM1(6332) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM1(6332))))  severity failure;
	assert RAM1(6333) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM1(6333))))  severity failure;
	assert RAM1(6334) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM1(6334))))  severity failure;
	assert RAM1(6335) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM1(6335))))  severity failure;
	assert RAM1(6336) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM1(6336))))  severity failure;
	assert RAM1(6337) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM1(6337))))  severity failure;
	assert RAM1(6338) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM1(6338))))  severity failure;
	assert RAM1(6339) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM1(6339))))  severity failure;
	assert RAM1(6340) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM1(6340))))  severity failure;
	assert RAM1(6341) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM1(6341))))  severity failure;
	assert RAM1(6342) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM1(6342))))  severity failure;
	assert RAM1(6343) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM1(6343))))  severity failure;
	assert RAM1(6344) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM1(6344))))  severity failure;
	assert RAM1(6345) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM1(6345))))  severity failure;
	assert RAM1(6346) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM1(6346))))  severity failure;
	assert RAM1(6347) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM1(6347))))  severity failure;
	assert RAM1(6348) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM1(6348))))  severity failure;
	assert RAM1(6349) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM1(6349))))  severity failure;
	assert RAM1(6350) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM1(6350))))  severity failure;
	assert RAM1(6351) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM1(6351))))  severity failure;
	assert RAM1(6352) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM1(6352))))  severity failure;
	assert RAM1(6353) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM1(6353))))  severity failure;
	assert RAM1(6354) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM1(6354))))  severity failure;
	assert RAM1(6355) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM1(6355))))  severity failure;
	assert RAM1(6356) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM1(6356))))  severity failure;
	assert RAM1(6357) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM1(6357))))  severity failure;
	assert RAM1(6358) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM1(6358))))  severity failure;
	assert RAM1(6359) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM1(6359))))  severity failure;
	assert RAM1(6360) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM1(6360))))  severity failure;
	assert RAM1(6361) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM1(6361))))  severity failure;
	assert RAM1(6362) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM1(6362))))  severity failure;
	assert RAM1(6363) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM1(6363))))  severity failure;
	assert RAM1(6364) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM1(6364))))  severity failure;
	assert RAM1(6365) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM1(6365))))  severity failure;
	assert RAM1(6366) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM1(6366))))  severity failure;
	assert RAM1(6367) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM1(6367))))  severity failure;
	assert RAM1(6368) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM1(6368))))  severity failure;
	assert RAM1(6369) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM1(6369))))  severity failure;
	assert RAM1(6370) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM1(6370))))  severity failure;
	assert RAM1(6371) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM1(6371))))  severity failure;
	assert RAM1(6372) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM1(6372))))  severity failure;
	assert RAM1(6373) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM1(6373))))  severity failure;
	assert RAM1(6374) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM1(6374))))  severity failure;
	assert RAM1(6375) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM1(6375))))  severity failure;
	assert RAM1(6376) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM1(6376))))  severity failure;
	assert RAM1(6377) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM1(6377))))  severity failure;
	assert RAM1(6378) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM1(6378))))  severity failure;
	assert RAM1(6379) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM1(6379))))  severity failure;
	assert RAM1(6380) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM1(6380))))  severity failure;
	assert RAM1(6381) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM1(6381))))  severity failure;
	assert RAM1(6382) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM1(6382))))  severity failure;
	assert RAM1(6383) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM1(6383))))  severity failure;
	assert RAM1(6384) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM1(6384))))  severity failure;
	assert RAM1(6385) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM1(6385))))  severity failure;
	assert RAM1(6386) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM1(6386))))  severity failure;
	assert RAM1(6387) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM1(6387))))  severity failure;
	assert RAM1(6388) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM1(6388))))  severity failure;
	assert RAM1(6389) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM1(6389))))  severity failure;
	assert RAM1(6390) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM1(6390))))  severity failure;
	assert RAM1(6391) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM1(6391))))  severity failure;
	assert RAM1(6392) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM1(6392))))  severity failure;
	assert RAM1(6393) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM1(6393))))  severity failure;
	assert RAM1(6394) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM1(6394))))  severity failure;
	assert RAM1(6395) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM1(6395))))  severity failure;
	assert RAM1(6396) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM1(6396))))  severity failure;
	assert RAM1(6397) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM1(6397))))  severity failure;
	assert RAM1(6398) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM1(6398))))  severity failure;
	assert RAM1(6399) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM1(6399))))  severity failure;
	assert RAM1(6400) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM1(6400))))  severity failure;
	assert RAM1(6401) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM1(6401))))  severity failure;
	assert RAM1(6402) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM1(6402))))  severity failure;
	assert RAM1(6403) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM1(6403))))  severity failure;
	assert RAM1(6404) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM1(6404))))  severity failure;
	assert RAM1(6405) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM1(6405))))  severity failure;
	assert RAM1(6406) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM1(6406))))  severity failure;
	assert RAM1(6407) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM1(6407))))  severity failure;
	assert RAM1(6408) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM1(6408))))  severity failure;
	assert RAM1(6409) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM1(6409))))  severity failure;
	assert RAM1(6410) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM1(6410))))  severity failure;
	assert RAM1(6411) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM1(6411))))  severity failure;
	assert RAM1(6412) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM1(6412))))  severity failure;
	assert RAM1(6413) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM1(6413))))  severity failure;
	assert RAM1(6414) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM1(6414))))  severity failure;
	assert RAM1(6415) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM1(6415))))  severity failure;
	assert RAM1(6416) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM1(6416))))  severity failure;
	assert RAM1(6417) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM1(6417))))  severity failure;
	assert RAM1(6418) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM1(6418))))  severity failure;
	assert RAM1(6419) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM1(6419))))  severity failure;
	assert RAM1(6420) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM1(6420))))  severity failure;
	assert RAM1(6421) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM1(6421))))  severity failure;
	assert RAM1(6422) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM1(6422))))  severity failure;
	assert RAM1(6423) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM1(6423))))  severity failure;
	assert RAM1(6424) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM1(6424))))  severity failure;
	assert RAM1(6425) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM1(6425))))  severity failure;
	assert RAM1(6426) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM1(6426))))  severity failure;
	assert RAM1(6427) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM1(6427))))  severity failure;
	assert RAM1(6428) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM1(6428))))  severity failure;
	assert RAM1(6429) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM1(6429))))  severity failure;
	assert RAM1(6430) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM1(6430))))  severity failure;
	assert RAM1(6431) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM1(6431))))  severity failure;
	assert RAM1(6432) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM1(6432))))  severity failure;
	assert RAM1(6433) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM1(6433))))  severity failure;
	assert RAM1(6434) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM1(6434))))  severity failure;
	assert RAM1(6435) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM1(6435))))  severity failure;
	assert RAM1(6436) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM1(6436))))  severity failure;
	assert RAM1(6437) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM1(6437))))  severity failure;
	assert RAM1(6438) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM1(6438))))  severity failure;
	assert RAM1(6439) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM1(6439))))  severity failure;
	assert RAM1(6440) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM1(6440))))  severity failure;
	assert RAM1(6441) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM1(6441))))  severity failure;
	assert RAM1(6442) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM1(6442))))  severity failure;
	assert RAM1(6443) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM1(6443))))  severity failure;
	assert RAM1(6444) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM1(6444))))  severity failure;
	assert RAM1(6445) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM1(6445))))  severity failure;
	assert RAM1(6446) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM1(6446))))  severity failure;
	assert RAM1(6447) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM1(6447))))  severity failure;
	assert RAM1(6448) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM1(6448))))  severity failure;
	assert RAM1(6449) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM1(6449))))  severity failure;
	assert RAM1(6450) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM1(6450))))  severity failure;
	assert RAM1(6451) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM1(6451))))  severity failure;
	assert RAM1(6452) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM1(6452))))  severity failure;
	assert RAM1(6453) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM1(6453))))  severity failure;
	assert RAM1(6454) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM1(6454))))  severity failure;
	assert RAM1(6455) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM1(6455))))  severity failure;
	assert RAM1(6456) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM1(6456))))  severity failure;
	assert RAM1(6457) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM1(6457))))  severity failure;
	assert RAM1(6458) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM1(6458))))  severity failure;
	assert RAM1(6459) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM1(6459))))  severity failure;
	assert RAM1(6460) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM1(6460))))  severity failure;
	assert RAM1(6461) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM1(6461))))  severity failure;
	assert RAM1(6462) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM1(6462))))  severity failure;
	assert RAM1(6463) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM1(6463))))  severity failure;
	assert RAM1(6464) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM1(6464))))  severity failure;
	assert RAM1(6465) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM1(6465))))  severity failure;
	assert RAM1(6466) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM1(6466))))  severity failure;
	assert RAM1(6467) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM1(6467))))  severity failure;
	assert RAM1(6468) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM1(6468))))  severity failure;
	assert RAM1(6469) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM1(6469))))  severity failure;
	assert RAM1(6470) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM1(6470))))  severity failure;
	assert RAM1(6471) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM1(6471))))  severity failure;
	assert RAM1(6472) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM1(6472))))  severity failure;
	assert RAM1(6473) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM1(6473))))  severity failure;
	assert RAM1(6474) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM1(6474))))  severity failure;
	assert RAM1(6475) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM1(6475))))  severity failure;
	assert RAM1(6476) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM1(6476))))  severity failure;
	assert RAM1(6477) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM1(6477))))  severity failure;
	assert RAM1(6478) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM1(6478))))  severity failure;
	assert RAM1(6479) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM1(6479))))  severity failure;
	assert RAM1(6480) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM1(6480))))  severity failure;
	assert RAM1(6481) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM1(6481))))  severity failure;
	assert RAM1(6482) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM1(6482))))  severity failure;
	assert RAM1(6483) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM1(6483))))  severity failure;
	assert RAM1(6484) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM1(6484))))  severity failure;
	assert RAM1(6485) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM1(6485))))  severity failure;
	assert RAM1(6486) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM1(6486))))  severity failure;
	assert RAM1(6487) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM1(6487))))  severity failure;
	assert RAM1(6488) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM1(6488))))  severity failure;
	assert RAM1(6489) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM1(6489))))  severity failure;
	assert RAM1(6490) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM1(6490))))  severity failure;
	assert RAM1(6491) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM1(6491))))  severity failure;
	assert RAM1(6492) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM1(6492))))  severity failure;
	assert RAM1(6493) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM1(6493))))  severity failure;
	assert RAM1(6494) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM1(6494))))  severity failure;
	assert RAM1(6495) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM1(6495))))  severity failure;
	assert RAM1(6496) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM1(6496))))  severity failure;
	assert RAM1(6497) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM1(6497))))  severity failure;
	assert RAM1(6498) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM1(6498))))  severity failure;
	assert RAM1(6499) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM1(6499))))  severity failure;
	assert RAM1(6500) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM1(6500))))  severity failure;
	assert RAM1(6501) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM1(6501))))  severity failure;
	assert RAM1(6502) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM1(6502))))  severity failure;
	assert RAM1(6503) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM1(6503))))  severity failure;
	assert RAM1(6504) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM1(6504))))  severity failure;
	assert RAM1(6505) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM1(6505))))  severity failure;
	assert RAM1(6506) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM1(6506))))  severity failure;
	assert RAM1(6507) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM1(6507))))  severity failure;
	assert RAM1(6508) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM1(6508))))  severity failure;
	assert RAM1(6509) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM1(6509))))  severity failure;
	assert RAM1(6510) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM1(6510))))  severity failure;
	assert RAM1(6511) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM1(6511))))  severity failure;
	assert RAM1(6512) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM1(6512))))  severity failure;
	assert RAM1(6513) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM1(6513))))  severity failure;
	assert RAM1(6514) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM1(6514))))  severity failure;
	assert RAM1(6515) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM1(6515))))  severity failure;
	assert RAM1(6516) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM1(6516))))  severity failure;
	assert RAM1(6517) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM1(6517))))  severity failure;
	assert RAM1(6518) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM1(6518))))  severity failure;
	assert RAM1(6519) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM1(6519))))  severity failure;
	assert RAM1(6520) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM1(6520))))  severity failure;
	assert RAM1(6521) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM1(6521))))  severity failure;
	assert RAM1(6522) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM1(6522))))  severity failure;
	assert RAM1(6523) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM1(6523))))  severity failure;
	assert RAM1(6524) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM1(6524))))  severity failure;
	assert RAM1(6525) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM1(6525))))  severity failure;
	assert RAM1(6526) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM1(6526))))  severity failure;
	assert RAM1(6527) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM1(6527))))  severity failure;
	assert RAM1(6528) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM1(6528))))  severity failure;
	assert RAM1(6529) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM1(6529))))  severity failure;
	assert RAM1(6530) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM1(6530))))  severity failure;
	assert RAM1(6531) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM1(6531))))  severity failure;
	assert RAM1(6532) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM1(6532))))  severity failure;
	assert RAM1(6533) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM1(6533))))  severity failure;
	assert RAM1(6534) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM1(6534))))  severity failure;
	assert RAM1(6535) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM1(6535))))  severity failure;
	assert RAM1(6536) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM1(6536))))  severity failure;
	assert RAM1(6537) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM1(6537))))  severity failure;
	assert RAM1(6538) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM1(6538))))  severity failure;
	assert RAM1(6539) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM1(6539))))  severity failure;
	assert RAM1(6540) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM1(6540))))  severity failure;
	assert RAM1(6541) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM1(6541))))  severity failure;
	assert RAM1(6542) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM1(6542))))  severity failure;
	assert RAM1(6543) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM1(6543))))  severity failure;
	assert RAM1(6544) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM1(6544))))  severity failure;
	assert RAM1(6545) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM1(6545))))  severity failure;
	assert RAM1(6546) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM1(6546))))  severity failure;
	assert RAM1(6547) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM1(6547))))  severity failure;
	assert RAM1(6548) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM1(6548))))  severity failure;
	assert RAM1(6549) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM1(6549))))  severity failure;
	assert RAM1(6550) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM1(6550))))  severity failure;
	assert RAM1(6551) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM1(6551))))  severity failure;
	assert RAM1(6552) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM1(6552))))  severity failure;
	assert RAM1(6553) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM1(6553))))  severity failure;
	assert RAM1(6554) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM1(6554))))  severity failure;
	assert RAM1(6555) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM1(6555))))  severity failure;
	assert RAM1(6556) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM1(6556))))  severity failure;
	assert RAM1(6557) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM1(6557))))  severity failure;
	assert RAM1(6558) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM1(6558))))  severity failure;
	assert RAM1(6559) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM1(6559))))  severity failure;
	assert RAM1(6560) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM1(6560))))  severity failure;
	assert RAM1(6561) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM1(6561))))  severity failure;
	assert RAM1(6562) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM1(6562))))  severity failure;
	assert RAM1(6563) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM1(6563))))  severity failure;
	assert RAM1(6564) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM1(6564))))  severity failure;
	assert RAM1(6565) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM1(6565))))  severity failure;
	assert RAM1(6566) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM1(6566))))  severity failure;
	assert RAM1(6567) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM1(6567))))  severity failure;
	assert RAM1(6568) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM1(6568))))  severity failure;
	assert RAM1(6569) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM1(6569))))  severity failure;
	assert RAM1(6570) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM1(6570))))  severity failure;
	assert RAM1(6571) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM1(6571))))  severity failure;
	assert RAM1(6572) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM1(6572))))  severity failure;
	assert RAM1(6573) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM1(6573))))  severity failure;
	assert RAM1(6574) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM1(6574))))  severity failure;
	assert RAM1(6575) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM1(6575))))  severity failure;
	assert RAM1(6576) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM1(6576))))  severity failure;
	assert RAM1(6577) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM1(6577))))  severity failure;
	assert RAM1(6578) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM1(6578))))  severity failure;
	assert RAM1(6579) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM1(6579))))  severity failure;
	assert RAM1(6580) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM1(6580))))  severity failure;
	assert RAM1(6581) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM1(6581))))  severity failure;
	assert RAM1(6582) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM1(6582))))  severity failure;
	assert RAM1(6583) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM1(6583))))  severity failure;
	assert RAM1(6584) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM1(6584))))  severity failure;
	assert RAM1(6585) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM1(6585))))  severity failure;
	assert RAM1(6586) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM1(6586))))  severity failure;
	assert RAM1(6587) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM1(6587))))  severity failure;
	assert RAM1(6588) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM1(6588))))  severity failure;
	assert RAM1(6589) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM1(6589))))  severity failure;
	assert RAM1(6590) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM1(6590))))  severity failure;
	assert RAM1(6591) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM1(6591))))  severity failure;
	assert RAM1(6592) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM1(6592))))  severity failure;
	assert RAM1(6593) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM1(6593))))  severity failure;
	assert RAM1(6594) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM1(6594))))  severity failure;
	assert RAM1(6595) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM1(6595))))  severity failure;
	assert RAM1(6596) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM1(6596))))  severity failure;
	assert RAM1(6597) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM1(6597))))  severity failure;
	assert RAM1(6598) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM1(6598))))  severity failure;
	assert RAM1(6599) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM1(6599))))  severity failure;
	assert RAM1(6600) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM1(6600))))  severity failure;
	assert RAM1(6601) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM1(6601))))  severity failure;
	assert RAM1(6602) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM1(6602))))  severity failure;
	assert RAM1(6603) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM1(6603))))  severity failure;
	assert RAM1(6604) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM1(6604))))  severity failure;
	assert RAM1(6605) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM1(6605))))  severity failure;
	assert RAM1(6606) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM1(6606))))  severity failure;
	assert RAM1(6607) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM1(6607))))  severity failure;
	assert RAM1(6608) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM1(6608))))  severity failure;
	assert RAM1(6609) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM1(6609))))  severity failure;
	assert RAM1(6610) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM1(6610))))  severity failure;
	assert RAM1(6611) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM1(6611))))  severity failure;
	assert RAM1(6612) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM1(6612))))  severity failure;
	assert RAM1(6613) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM1(6613))))  severity failure;
	assert RAM1(6614) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM1(6614))))  severity failure;
	assert RAM1(6615) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM1(6615))))  severity failure;
	assert RAM1(6616) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM1(6616))))  severity failure;
	assert RAM1(6617) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM1(6617))))  severity failure;
	assert RAM1(6618) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM1(6618))))  severity failure;
	assert RAM1(6619) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM1(6619))))  severity failure;
	assert RAM1(6620) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM1(6620))))  severity failure;
	assert RAM1(6621) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM1(6621))))  severity failure;
	assert RAM1(6622) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM1(6622))))  severity failure;
	assert RAM1(6623) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM1(6623))))  severity failure;
	assert RAM1(6624) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM1(6624))))  severity failure;
	assert RAM1(6625) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM1(6625))))  severity failure;
	assert RAM1(6626) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM1(6626))))  severity failure;
	assert RAM1(6627) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM1(6627))))  severity failure;
	assert RAM1(6628) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM1(6628))))  severity failure;
	assert RAM1(6629) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM1(6629))))  severity failure;
	assert RAM1(6630) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM1(6630))))  severity failure;
	assert RAM1(6631) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM1(6631))))  severity failure;
	assert RAM1(6632) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM1(6632))))  severity failure;
	assert RAM1(6633) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM1(6633))))  severity failure;
	assert RAM1(6634) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM1(6634))))  severity failure;
	assert RAM1(6635) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM1(6635))))  severity failure;
	assert RAM1(6636) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM1(6636))))  severity failure;
	assert RAM1(6637) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM1(6637))))  severity failure;
	assert RAM1(6638) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM1(6638))))  severity failure;
	assert RAM1(6639) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM1(6639))))  severity failure;
	assert RAM1(6640) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM1(6640))))  severity failure;
	assert RAM1(6641) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM1(6641))))  severity failure;
	assert RAM1(6642) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM1(6642))))  severity failure;
	assert RAM1(6643) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM1(6643))))  severity failure;
	assert RAM1(6644) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM1(6644))))  severity failure;
	assert RAM1(6645) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM1(6645))))  severity failure;
	assert RAM1(6646) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM1(6646))))  severity failure;
	assert RAM1(6647) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM1(6647))))  severity failure;
	assert RAM1(6648) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM1(6648))))  severity failure;
	assert RAM1(6649) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM1(6649))))  severity failure;
	assert RAM1(6650) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM1(6650))))  severity failure;
	assert RAM1(6651) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM1(6651))))  severity failure;
	assert RAM1(6652) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM1(6652))))  severity failure;
	assert RAM1(6653) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM1(6653))))  severity failure;
	assert RAM1(6654) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM1(6654))))  severity failure;
	assert RAM1(6655) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM1(6655))))  severity failure;
	assert RAM1(6656) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM1(6656))))  severity failure;
	assert RAM1(6657) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM1(6657))))  severity failure;
	assert RAM1(6658) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM1(6658))))  severity failure;
	assert RAM1(6659) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM1(6659))))  severity failure;
	assert RAM1(6660) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM1(6660))))  severity failure;
	assert RAM1(6661) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM1(6661))))  severity failure;
	assert RAM1(6662) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM1(6662))))  severity failure;
	assert RAM1(6663) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM1(6663))))  severity failure;
	assert RAM1(6664) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM1(6664))))  severity failure;
	assert RAM1(6665) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM1(6665))))  severity failure;
	assert RAM1(6666) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM1(6666))))  severity failure;
	assert RAM1(6667) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM1(6667))))  severity failure;
	assert RAM1(6668) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM1(6668))))  severity failure;
	assert RAM1(6669) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM1(6669))))  severity failure;
	assert RAM1(6670) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM1(6670))))  severity failure;
	assert RAM1(6671) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM1(6671))))  severity failure;
	assert RAM1(6672) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM1(6672))))  severity failure;
	assert RAM1(6673) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM1(6673))))  severity failure;
	assert RAM1(6674) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM1(6674))))  severity failure;
	assert RAM1(6675) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM1(6675))))  severity failure;
	assert RAM1(6676) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM1(6676))))  severity failure;
	assert RAM1(6677) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM1(6677))))  severity failure;
	assert RAM1(6678) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM1(6678))))  severity failure;
	assert RAM1(6679) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM1(6679))))  severity failure;
	assert RAM1(6680) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM1(6680))))  severity failure;
	assert RAM1(6681) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM1(6681))))  severity failure;
	assert RAM1(6682) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM1(6682))))  severity failure;
	assert RAM1(6683) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM1(6683))))  severity failure;
	assert RAM1(6684) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM1(6684))))  severity failure;
	assert RAM1(6685) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM1(6685))))  severity failure;
	assert RAM1(6686) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM1(6686))))  severity failure;
	assert RAM1(6687) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM1(6687))))  severity failure;
	assert RAM1(6688) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM1(6688))))  severity failure;
	assert RAM1(6689) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM1(6689))))  severity failure;
	assert RAM1(6690) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM1(6690))))  severity failure;
	assert RAM1(6691) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM1(6691))))  severity failure;
	assert RAM1(6692) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM1(6692))))  severity failure;
	assert RAM1(6693) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM1(6693))))  severity failure;
	assert RAM1(6694) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM1(6694))))  severity failure;
	assert RAM1(6695) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM1(6695))))  severity failure;
	assert RAM1(6696) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM1(6696))))  severity failure;
	assert RAM1(6697) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM1(6697))))  severity failure;
	assert RAM1(6698) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM1(6698))))  severity failure;
	assert RAM1(6699) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM1(6699))))  severity failure;
	assert RAM1(6700) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM1(6700))))  severity failure;
	assert RAM1(6701) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM1(6701))))  severity failure;
	assert RAM1(6702) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM1(6702))))  severity failure;
	assert RAM1(6703) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM1(6703))))  severity failure;
	assert RAM1(6704) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM1(6704))))  severity failure;
	assert RAM1(6705) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM1(6705))))  severity failure;
	assert RAM1(6706) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM1(6706))))  severity failure;
	assert RAM1(6707) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM1(6707))))  severity failure;
	assert RAM1(6708) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM1(6708))))  severity failure;
	assert RAM1(6709) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM1(6709))))  severity failure;
	assert RAM1(6710) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM1(6710))))  severity failure;
	assert RAM1(6711) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM1(6711))))  severity failure;
	assert RAM1(6712) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM1(6712))))  severity failure;
	assert RAM1(6713) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM1(6713))))  severity failure;
	assert RAM1(6714) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM1(6714))))  severity failure;
	assert RAM1(6715) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM1(6715))))  severity failure;
	assert RAM1(6716) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM1(6716))))  severity failure;
	assert RAM1(6717) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM1(6717))))  severity failure;
	assert RAM1(6718) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM1(6718))))  severity failure;
	assert RAM1(6719) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM1(6719))))  severity failure;
	assert RAM1(6720) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM1(6720))))  severity failure;
	assert RAM1(6721) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM1(6721))))  severity failure;
	assert RAM1(6722) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM1(6722))))  severity failure;
	assert RAM1(6723) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM1(6723))))  severity failure;
	assert RAM1(6724) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM1(6724))))  severity failure;
	assert RAM1(6725) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM1(6725))))  severity failure;
	assert RAM1(6726) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM1(6726))))  severity failure;
	assert RAM1(6727) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM1(6727))))  severity failure;
	assert RAM1(6728) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM1(6728))))  severity failure;
	assert RAM1(6729) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM1(6729))))  severity failure;
	assert RAM1(6730) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM1(6730))))  severity failure;
	assert RAM1(6731) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM1(6731))))  severity failure;
	assert RAM1(6732) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM1(6732))))  severity failure;
	assert RAM1(6733) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM1(6733))))  severity failure;
	assert RAM1(6734) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM1(6734))))  severity failure;
	assert RAM1(6735) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM1(6735))))  severity failure;
	assert RAM1(6736) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM1(6736))))  severity failure;
	assert RAM1(6737) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM1(6737))))  severity failure;
	assert RAM1(6738) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM1(6738))))  severity failure;
	assert RAM1(6739) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM1(6739))))  severity failure;
	assert RAM1(6740) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM1(6740))))  severity failure;
	assert RAM1(6741) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM1(6741))))  severity failure;
	assert RAM1(6742) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM1(6742))))  severity failure;
	assert RAM1(6743) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM1(6743))))  severity failure;
	assert RAM1(6744) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM1(6744))))  severity failure;
	assert RAM1(6745) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM1(6745))))  severity failure;
	assert RAM1(6746) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM1(6746))))  severity failure;
	assert RAM1(6747) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM1(6747))))  severity failure;
	assert RAM1(6748) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM1(6748))))  severity failure;
	assert RAM1(6749) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM1(6749))))  severity failure;
	assert RAM1(6750) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM1(6750))))  severity failure;
	assert RAM1(6751) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM1(6751))))  severity failure;
	assert RAM1(6752) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM1(6752))))  severity failure;
	assert RAM1(6753) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM1(6753))))  severity failure;
	assert RAM1(6754) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM1(6754))))  severity failure;
	assert RAM1(6755) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM1(6755))))  severity failure;
	assert RAM1(6756) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM1(6756))))  severity failure;
	assert RAM1(6757) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM1(6757))))  severity failure;
	assert RAM1(6758) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM1(6758))))  severity failure;
	assert RAM1(6759) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM1(6759))))  severity failure;
	assert RAM1(6760) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM1(6760))))  severity failure;
	assert RAM1(6761) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM1(6761))))  severity failure;
	assert RAM1(6762) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM1(6762))))  severity failure;
	assert RAM1(6763) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM1(6763))))  severity failure;
	assert RAM1(6764) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM1(6764))))  severity failure;
	assert RAM1(6765) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM1(6765))))  severity failure;
	assert RAM1(6766) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM1(6766))))  severity failure;
	assert RAM1(6767) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM1(6767))))  severity failure;
	assert RAM1(6768) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM1(6768))))  severity failure;
	assert RAM1(6769) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM1(6769))))  severity failure;
	assert RAM1(6770) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM1(6770))))  severity failure;
	assert RAM1(6771) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM1(6771))))  severity failure;
	assert RAM1(6772) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM1(6772))))  severity failure;
	assert RAM1(6773) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM1(6773))))  severity failure;
	assert RAM1(6774) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM1(6774))))  severity failure;
	assert RAM1(6775) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM1(6775))))  severity failure;
	assert RAM1(6776) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM1(6776))))  severity failure;
	assert RAM1(6777) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM1(6777))))  severity failure;
	assert RAM1(6778) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM1(6778))))  severity failure;
	assert RAM1(6779) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM1(6779))))  severity failure;
	assert RAM1(6780) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM1(6780))))  severity failure;
	assert RAM1(6781) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM1(6781))))  severity failure;
	assert RAM1(6782) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM1(6782))))  severity failure;
	assert RAM1(6783) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM1(6783))))  severity failure;
	assert RAM1(6784) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM1(6784))))  severity failure;
	assert RAM1(6785) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM1(6785))))  severity failure;
	assert RAM1(6786) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM1(6786))))  severity failure;
	assert RAM1(6787) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM1(6787))))  severity failure;
	assert RAM1(6788) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM1(6788))))  severity failure;
	assert RAM1(6789) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM1(6789))))  severity failure;
	assert RAM1(6790) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM1(6790))))  severity failure;
	assert RAM1(6791) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM1(6791))))  severity failure;
	assert RAM1(6792) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM1(6792))))  severity failure;
	assert RAM1(6793) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM1(6793))))  severity failure;
	assert RAM1(6794) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM1(6794))))  severity failure;
	assert RAM1(6795) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM1(6795))))  severity failure;
	assert RAM1(6796) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM1(6796))))  severity failure;
	assert RAM1(6797) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM1(6797))))  severity failure;
	assert RAM1(6798) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM1(6798))))  severity failure;
	assert RAM1(6799) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM1(6799))))  severity failure;
	assert RAM1(6800) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM1(6800))))  severity failure;
	assert RAM1(6801) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM1(6801))))  severity failure;
	assert RAM1(6802) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM1(6802))))  severity failure;
	assert RAM1(6803) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM1(6803))))  severity failure;
	assert RAM1(6804) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM1(6804))))  severity failure;
	assert RAM1(6805) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM1(6805))))  severity failure;
	assert RAM1(6806) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM1(6806))))  severity failure;
	assert RAM1(6807) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM1(6807))))  severity failure;
	assert RAM1(6808) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM1(6808))))  severity failure;
	assert RAM1(6809) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM1(6809))))  severity failure;
	assert RAM1(6810) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM1(6810))))  severity failure;
	assert RAM1(6811) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM1(6811))))  severity failure;
	assert RAM1(6812) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM1(6812))))  severity failure;
	assert RAM1(6813) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM1(6813))))  severity failure;
	assert RAM1(6814) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM1(6814))))  severity failure;
	assert RAM1(6815) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM1(6815))))  severity failure;
	assert RAM1(6816) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM1(6816))))  severity failure;
	assert RAM1(6817) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM1(6817))))  severity failure;
	assert RAM1(6818) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM1(6818))))  severity failure;
	assert RAM1(6819) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM1(6819))))  severity failure;
	assert RAM1(6820) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM1(6820))))  severity failure;
	assert RAM1(6821) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM1(6821))))  severity failure;
	assert RAM1(6822) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM1(6822))))  severity failure;
	assert RAM1(6823) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM1(6823))))  severity failure;
	assert RAM1(6824) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM1(6824))))  severity failure;
	assert RAM1(6825) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM1(6825))))  severity failure;
	assert RAM1(6826) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM1(6826))))  severity failure;
	assert RAM1(6827) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM1(6827))))  severity failure;
	assert RAM1(6828) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM1(6828))))  severity failure;
	assert RAM1(6829) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM1(6829))))  severity failure;
	assert RAM1(6830) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM1(6830))))  severity failure;
	assert RAM1(6831) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM1(6831))))  severity failure;
	assert RAM1(6832) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM1(6832))))  severity failure;
	assert RAM1(6833) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM1(6833))))  severity failure;
	assert RAM1(6834) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM1(6834))))  severity failure;
	assert RAM1(6835) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM1(6835))))  severity failure;
	assert RAM1(6836) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM1(6836))))  severity failure;
	assert RAM1(6837) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM1(6837))))  severity failure;
	assert RAM1(6838) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM1(6838))))  severity failure;
	assert RAM1(6839) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM1(6839))))  severity failure;
	assert RAM1(6840) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM1(6840))))  severity failure;
	assert RAM1(6841) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM1(6841))))  severity failure;
	assert RAM1(6842) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM1(6842))))  severity failure;
	assert RAM1(6843) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM1(6843))))  severity failure;
	assert RAM1(6844) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM1(6844))))  severity failure;
	assert RAM1(6845) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM1(6845))))  severity failure;
	assert RAM1(6846) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM1(6846))))  severity failure;
	assert RAM1(6847) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM1(6847))))  severity failure;
	assert RAM1(6848) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM1(6848))))  severity failure;
	assert RAM1(6849) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM1(6849))))  severity failure;
	assert RAM1(6850) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM1(6850))))  severity failure;
	assert RAM1(6851) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM1(6851))))  severity failure;
	assert RAM1(6852) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM1(6852))))  severity failure;
	assert RAM1(6853) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM1(6853))))  severity failure;
	assert RAM1(6854) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM1(6854))))  severity failure;
	assert RAM1(6855) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM1(6855))))  severity failure;
	assert RAM1(6856) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM1(6856))))  severity failure;
	assert RAM1(6857) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM1(6857))))  severity failure;
	assert RAM1(6858) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM1(6858))))  severity failure;
	assert RAM1(6859) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM1(6859))))  severity failure;
	assert RAM1(6860) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM1(6860))))  severity failure;
	assert RAM1(6861) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM1(6861))))  severity failure;
	assert RAM1(6862) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM1(6862))))  severity failure;
	assert RAM1(6863) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM1(6863))))  severity failure;
	assert RAM1(6864) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM1(6864))))  severity failure;
	assert RAM1(6865) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM1(6865))))  severity failure;
	assert RAM1(6866) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM1(6866))))  severity failure;
	assert RAM1(6867) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM1(6867))))  severity failure;
	assert RAM1(6868) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM1(6868))))  severity failure;
	assert RAM1(6869) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM1(6869))))  severity failure;
	assert RAM1(6870) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM1(6870))))  severity failure;
	assert RAM1(6871) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM1(6871))))  severity failure;
	assert RAM1(6872) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM1(6872))))  severity failure;
	assert RAM1(6873) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM1(6873))))  severity failure;
	assert RAM1(6874) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM1(6874))))  severity failure;
	assert RAM1(6875) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM1(6875))))  severity failure;
	assert RAM1(6876) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM1(6876))))  severity failure;
	assert RAM1(6877) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM1(6877))))  severity failure;
	assert RAM1(6878) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM1(6878))))  severity failure;
	assert RAM1(6879) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM1(6879))))  severity failure;
	assert RAM1(6880) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM1(6880))))  severity failure;
	assert RAM1(6881) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM1(6881))))  severity failure;
	assert RAM1(6882) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM1(6882))))  severity failure;
	assert RAM1(6883) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM1(6883))))  severity failure;
	assert RAM1(6884) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM1(6884))))  severity failure;
	assert RAM1(6885) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM1(6885))))  severity failure;
	assert RAM1(6886) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM1(6886))))  severity failure;
	assert RAM1(6887) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM1(6887))))  severity failure;
	assert RAM1(6888) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM1(6888))))  severity failure;
	assert RAM1(6889) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM1(6889))))  severity failure;
	assert RAM1(6890) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM1(6890))))  severity failure;
	assert RAM1(6891) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM1(6891))))  severity failure;
	assert RAM1(6892) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM1(6892))))  severity failure;
	assert RAM1(6893) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM1(6893))))  severity failure;
	assert RAM1(6894) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM1(6894))))  severity failure;
	assert RAM1(6895) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM1(6895))))  severity failure;
	assert RAM1(6896) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM1(6896))))  severity failure;
	assert RAM1(6897) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM1(6897))))  severity failure;
	assert RAM1(6898) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM1(6898))))  severity failure;
	assert RAM1(6899) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM1(6899))))  severity failure;
	assert RAM1(6900) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM1(6900))))  severity failure;
	assert RAM1(6901) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM1(6901))))  severity failure;
	assert RAM1(6902) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM1(6902))))  severity failure;
	assert RAM1(6903) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM1(6903))))  severity failure;
	assert RAM1(6904) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM1(6904))))  severity failure;
	assert RAM1(6905) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM1(6905))))  severity failure;
	assert RAM1(6906) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM1(6906))))  severity failure;
	assert RAM1(6907) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM1(6907))))  severity failure;
	assert RAM1(6908) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM1(6908))))  severity failure;
	assert RAM1(6909) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM1(6909))))  severity failure;
	assert RAM1(6910) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM1(6910))))  severity failure;
	assert RAM1(6911) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM1(6911))))  severity failure;
	assert RAM1(6912) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM1(6912))))  severity failure;
	assert RAM1(6913) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM1(6913))))  severity failure;
	assert RAM1(6914) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM1(6914))))  severity failure;
	assert RAM1(6915) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM1(6915))))  severity failure;
	assert RAM1(6916) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM1(6916))))  severity failure;
	assert RAM1(6917) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM1(6917))))  severity failure;
	assert RAM1(6918) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM1(6918))))  severity failure;
	assert RAM1(6919) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM1(6919))))  severity failure;
	assert RAM1(6920) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM1(6920))))  severity failure;
	assert RAM1(6921) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM1(6921))))  severity failure;
	assert RAM1(6922) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM1(6922))))  severity failure;
	assert RAM1(6923) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM1(6923))))  severity failure;
	assert RAM1(6924) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM1(6924))))  severity failure;
	assert RAM1(6925) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM1(6925))))  severity failure;
	assert RAM1(6926) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM1(6926))))  severity failure;
	assert RAM1(6927) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM1(6927))))  severity failure;
	assert RAM1(6928) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM1(6928))))  severity failure;
	assert RAM1(6929) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM1(6929))))  severity failure;
	assert RAM1(6930) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM1(6930))))  severity failure;
	assert RAM1(6931) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM1(6931))))  severity failure;
	assert RAM1(6932) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM1(6932))))  severity failure;
	assert RAM1(6933) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM1(6933))))  severity failure;
	assert RAM1(6934) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM1(6934))))  severity failure;
	assert RAM1(6935) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM1(6935))))  severity failure;
	assert RAM1(6936) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM1(6936))))  severity failure;
	assert RAM1(6937) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM1(6937))))  severity failure;
	assert RAM1(6938) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM1(6938))))  severity failure;
	assert RAM1(6939) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM1(6939))))  severity failure;
	assert RAM1(6940) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM1(6940))))  severity failure;
	assert RAM1(6941) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM1(6941))))  severity failure;
	assert RAM1(6942) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM1(6942))))  severity failure;
	assert RAM1(6943) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM1(6943))))  severity failure;
	assert RAM1(6944) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM1(6944))))  severity failure;
	assert RAM1(6945) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM1(6945))))  severity failure;
	assert RAM1(6946) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM1(6946))))  severity failure;
	assert RAM1(6947) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM1(6947))))  severity failure;
	assert RAM1(6948) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM1(6948))))  severity failure;
	assert RAM1(6949) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM1(6949))))  severity failure;
	assert RAM1(6950) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM1(6950))))  severity failure;
	assert RAM1(6951) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM1(6951))))  severity failure;
	assert RAM1(6952) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM1(6952))))  severity failure;
	assert RAM1(6953) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM1(6953))))  severity failure;
	assert RAM1(6954) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM1(6954))))  severity failure;
	assert RAM1(6955) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM1(6955))))  severity failure;
	assert RAM1(6956) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM1(6956))))  severity failure;
	assert RAM1(6957) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM1(6957))))  severity failure;
	assert RAM1(6958) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM1(6958))))  severity failure;
	assert RAM1(6959) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM1(6959))))  severity failure;
	assert RAM1(6960) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM1(6960))))  severity failure;
	assert RAM1(6961) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM1(6961))))  severity failure;
	assert RAM1(6962) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM1(6962))))  severity failure;
	assert RAM1(6963) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM1(6963))))  severity failure;
	assert RAM1(6964) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM1(6964))))  severity failure;
	assert RAM1(6965) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM1(6965))))  severity failure;
	assert RAM1(6966) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM1(6966))))  severity failure;
	assert RAM1(6967) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM1(6967))))  severity failure;
	assert RAM1(6968) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM1(6968))))  severity failure;
	assert RAM1(6969) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM1(6969))))  severity failure;
	assert RAM1(6970) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM1(6970))))  severity failure;
	assert RAM1(6971) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM1(6971))))  severity failure;
	assert RAM1(6972) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM1(6972))))  severity failure;
	assert RAM1(6973) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM1(6973))))  severity failure;
	assert RAM1(6974) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM1(6974))))  severity failure;
	assert RAM1(6975) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM1(6975))))  severity failure;
	assert RAM1(6976) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM1(6976))))  severity failure;
	assert RAM1(6977) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM1(6977))))  severity failure;
	assert RAM1(6978) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM1(6978))))  severity failure;
	assert RAM1(6979) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM1(6979))))  severity failure;
	assert RAM1(6980) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM1(6980))))  severity failure;
	assert RAM1(6981) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM1(6981))))  severity failure;
	assert RAM1(6982) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM1(6982))))  severity failure;
	assert RAM1(6983) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM1(6983))))  severity failure;
	assert RAM1(6984) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM1(6984))))  severity failure;
	assert RAM1(6985) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM1(6985))))  severity failure;
	assert RAM1(6986) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM1(6986))))  severity failure;
	assert RAM1(6987) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM1(6987))))  severity failure;
	assert RAM1(6988) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM1(6988))))  severity failure;
	assert RAM1(6989) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM1(6989))))  severity failure;
	assert RAM1(6990) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM1(6990))))  severity failure;
	assert RAM1(6991) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM1(6991))))  severity failure;
	assert RAM1(6992) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM1(6992))))  severity failure;
	assert RAM1(6993) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM1(6993))))  severity failure;
	assert RAM1(6994) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM1(6994))))  severity failure;
	assert RAM1(6995) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM1(6995))))  severity failure;
	assert RAM1(6996) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM1(6996))))  severity failure;
	assert RAM1(6997) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM1(6997))))  severity failure;
	assert RAM1(6998) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM1(6998))))  severity failure;
	assert RAM1(6999) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM1(6999))))  severity failure;
	assert RAM1(7000) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM1(7000))))  severity failure;
	assert RAM1(7001) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM1(7001))))  severity failure;
	assert RAM1(7002) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM1(7002))))  severity failure;
	assert RAM1(7003) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM1(7003))))  severity failure;
	assert RAM1(7004) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM1(7004))))  severity failure;
	assert RAM1(7005) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM1(7005))))  severity failure;
	assert RAM1(7006) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM1(7006))))  severity failure;
	assert RAM1(7007) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM1(7007))))  severity failure;
	assert RAM1(7008) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM1(7008))))  severity failure;
	assert RAM1(7009) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM1(7009))))  severity failure;
	assert RAM1(7010) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM1(7010))))  severity failure;
	assert RAM1(7011) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM1(7011))))  severity failure;
	assert RAM1(7012) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM1(7012))))  severity failure;
	assert RAM1(7013) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM1(7013))))  severity failure;
	assert RAM1(7014) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM1(7014))))  severity failure;
	assert RAM1(7015) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM1(7015))))  severity failure;
	assert RAM1(7016) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM1(7016))))  severity failure;
	assert RAM1(7017) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM1(7017))))  severity failure;
	assert RAM1(7018) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM1(7018))))  severity failure;
	assert RAM1(7019) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM1(7019))))  severity failure;
	assert RAM1(7020) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM1(7020))))  severity failure;
	assert RAM1(7021) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM1(7021))))  severity failure;
	assert RAM1(7022) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM1(7022))))  severity failure;
	assert RAM1(7023) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM1(7023))))  severity failure;
	assert RAM1(7024) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM1(7024))))  severity failure;
	assert RAM1(7025) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM1(7025))))  severity failure;
	assert RAM1(7026) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM1(7026))))  severity failure;
	assert RAM1(7027) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM1(7027))))  severity failure;
	assert RAM1(7028) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM1(7028))))  severity failure;
	assert RAM1(7029) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM1(7029))))  severity failure;
	assert RAM1(7030) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM1(7030))))  severity failure;
	assert RAM1(7031) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM1(7031))))  severity failure;
	assert RAM1(7032) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM1(7032))))  severity failure;
	assert RAM1(7033) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM1(7033))))  severity failure;
	assert RAM1(7034) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM1(7034))))  severity failure;
	assert RAM1(7035) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM1(7035))))  severity failure;
	assert RAM1(7036) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM1(7036))))  severity failure;
	assert RAM1(7037) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM1(7037))))  severity failure;
	assert RAM1(7038) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM1(7038))))  severity failure;
	assert RAM1(7039) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM1(7039))))  severity failure;
	assert RAM1(7040) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM1(7040))))  severity failure;
	assert RAM1(7041) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM1(7041))))  severity failure;
	assert RAM1(7042) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM1(7042))))  severity failure;
	assert RAM1(7043) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM1(7043))))  severity failure;
	assert RAM1(7044) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM1(7044))))  severity failure;
	assert RAM1(7045) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM1(7045))))  severity failure;
	assert RAM1(7046) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM1(7046))))  severity failure;
	assert RAM1(7047) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM1(7047))))  severity failure;
	assert RAM1(7048) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM1(7048))))  severity failure;
	assert RAM1(7049) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM1(7049))))  severity failure;
	assert RAM1(7050) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM1(7050))))  severity failure;
	assert RAM1(7051) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM1(7051))))  severity failure;
	assert RAM1(7052) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM1(7052))))  severity failure;
	assert RAM1(7053) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM1(7053))))  severity failure;
	assert RAM1(7054) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM1(7054))))  severity failure;
	assert RAM1(7055) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM1(7055))))  severity failure;
	assert RAM1(7056) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM1(7056))))  severity failure;
	assert RAM1(7057) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM1(7057))))  severity failure;
	assert RAM1(7058) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM1(7058))))  severity failure;
	assert RAM1(7059) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM1(7059))))  severity failure;
	assert RAM1(7060) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM1(7060))))  severity failure;
	assert RAM1(7061) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM1(7061))))  severity failure;
	assert RAM1(7062) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM1(7062))))  severity failure;
	assert RAM1(7063) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM1(7063))))  severity failure;
	assert RAM1(7064) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM1(7064))))  severity failure;
	assert RAM1(7065) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM1(7065))))  severity failure;
	assert RAM1(7066) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM1(7066))))  severity failure;
	assert RAM1(7067) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM1(7067))))  severity failure;
	assert RAM1(7068) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM1(7068))))  severity failure;
	assert RAM1(7069) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM1(7069))))  severity failure;
	assert RAM1(7070) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM1(7070))))  severity failure;
	assert RAM1(7071) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM1(7071))))  severity failure;
	assert RAM1(7072) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM1(7072))))  severity failure;
	assert RAM1(7073) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM1(7073))))  severity failure;
	assert RAM1(7074) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM1(7074))))  severity failure;
	assert RAM1(7075) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM1(7075))))  severity failure;
	assert RAM1(7076) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM1(7076))))  severity failure;
	assert RAM1(7077) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM1(7077))))  severity failure;
	assert RAM1(7078) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM1(7078))))  severity failure;
	assert RAM1(7079) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM1(7079))))  severity failure;
	assert RAM1(7080) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM1(7080))))  severity failure;
	assert RAM1(7081) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM1(7081))))  severity failure;
	assert RAM1(7082) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM1(7082))))  severity failure;
	assert RAM1(7083) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM1(7083))))  severity failure;
	assert RAM1(7084) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM1(7084))))  severity failure;
	assert RAM1(7085) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM1(7085))))  severity failure;
	assert RAM1(7086) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM1(7086))))  severity failure;
	assert RAM1(7087) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM1(7087))))  severity failure;
	assert RAM1(7088) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM1(7088))))  severity failure;
	assert RAM1(7089) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM1(7089))))  severity failure;
	assert RAM1(7090) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM1(7090))))  severity failure;
	assert RAM1(7091) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM1(7091))))  severity failure;
	assert RAM1(7092) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM1(7092))))  severity failure;
	assert RAM1(7093) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM1(7093))))  severity failure;
	assert RAM1(7094) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM1(7094))))  severity failure;
	assert RAM1(7095) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM1(7095))))  severity failure;
	assert RAM1(7096) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM1(7096))))  severity failure;
	assert RAM1(7097) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM1(7097))))  severity failure;
	assert RAM1(7098) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM1(7098))))  severity failure;
	assert RAM1(7099) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM1(7099))))  severity failure;
	assert RAM1(7100) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM1(7100))))  severity failure;
	assert RAM1(7101) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM1(7101))))  severity failure;
	assert RAM1(7102) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM1(7102))))  severity failure;
	assert RAM1(7103) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM1(7103))))  severity failure;
	assert RAM1(7104) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM1(7104))))  severity failure;
	assert RAM1(7105) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM1(7105))))  severity failure;
	assert RAM1(7106) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM1(7106))))  severity failure;
	assert RAM1(7107) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM1(7107))))  severity failure;
	assert RAM1(7108) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM1(7108))))  severity failure;
	assert RAM1(7109) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM1(7109))))  severity failure;
	assert RAM1(7110) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM1(7110))))  severity failure;
	assert RAM1(7111) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM1(7111))))  severity failure;
	assert RAM1(7112) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM1(7112))))  severity failure;
	assert RAM1(7113) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM1(7113))))  severity failure;
	assert RAM1(7114) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM1(7114))))  severity failure;
	assert RAM1(7115) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM1(7115))))  severity failure;
	assert RAM1(7116) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM1(7116))))  severity failure;
	assert RAM1(7117) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM1(7117))))  severity failure;
	assert RAM1(7118) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM1(7118))))  severity failure;
	assert RAM1(7119) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM1(7119))))  severity failure;
	assert RAM1(7120) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM1(7120))))  severity failure;
	assert RAM1(7121) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM1(7121))))  severity failure;
	assert RAM1(7122) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM1(7122))))  severity failure;
	assert RAM1(7123) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM1(7123))))  severity failure;
	assert RAM1(7124) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM1(7124))))  severity failure;
	assert RAM1(7125) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM1(7125))))  severity failure;
	assert RAM1(7126) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM1(7126))))  severity failure;
	assert RAM1(7127) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM1(7127))))  severity failure;
	assert RAM1(7128) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM1(7128))))  severity failure;
	assert RAM1(7129) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM1(7129))))  severity failure;
	assert RAM1(7130) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM1(7130))))  severity failure;
	assert RAM1(7131) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM1(7131))))  severity failure;
	assert RAM1(7132) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM1(7132))))  severity failure;
	assert RAM1(7133) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM1(7133))))  severity failure;
	assert RAM1(7134) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM1(7134))))  severity failure;
	assert RAM1(7135) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM1(7135))))  severity failure;
	assert RAM1(7136) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM1(7136))))  severity failure;
	assert RAM1(7137) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM1(7137))))  severity failure;
	assert RAM1(7138) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM1(7138))))  severity failure;
	assert RAM1(7139) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM1(7139))))  severity failure;
	assert RAM1(7140) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM1(7140))))  severity failure;
	assert RAM1(7141) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM1(7141))))  severity failure;
	assert RAM1(7142) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM1(7142))))  severity failure;
	assert RAM1(7143) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM1(7143))))  severity failure;
	assert RAM1(7144) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM1(7144))))  severity failure;
	assert RAM1(7145) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM1(7145))))  severity failure;
	assert RAM1(7146) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM1(7146))))  severity failure;
	assert RAM1(7147) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM1(7147))))  severity failure;
	assert RAM1(7148) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM1(7148))))  severity failure;
	assert RAM1(7149) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM1(7149))))  severity failure;
	assert RAM1(7150) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM1(7150))))  severity failure;
	assert RAM1(7151) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM1(7151))))  severity failure;
	assert RAM1(7152) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM1(7152))))  severity failure;
	assert RAM1(7153) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM1(7153))))  severity failure;
	assert RAM1(7154) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM1(7154))))  severity failure;
	assert RAM1(7155) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM1(7155))))  severity failure;
	assert RAM1(7156) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM1(7156))))  severity failure;
	assert RAM1(7157) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM1(7157))))  severity failure;
	assert RAM1(7158) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM1(7158))))  severity failure;
	assert RAM1(7159) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM1(7159))))  severity failure;
	assert RAM1(7160) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM1(7160))))  severity failure;
	assert RAM1(7161) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM1(7161))))  severity failure;
	assert RAM1(7162) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM1(7162))))  severity failure;
	assert RAM1(7163) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM1(7163))))  severity failure;
	assert RAM1(7164) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM1(7164))))  severity failure;
	assert RAM1(7165) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM1(7165))))  severity failure;
	assert RAM1(7166) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM1(7166))))  severity failure;
	assert RAM1(7167) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM1(7167))))  severity failure;
	assert RAM1(7168) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM1(7168))))  severity failure;
	assert RAM1(7169) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM1(7169))))  severity failure;
	assert RAM1(7170) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM1(7170))))  severity failure;
	assert RAM1(7171) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM1(7171))))  severity failure;
	assert RAM1(7172) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM1(7172))))  severity failure;
	assert RAM1(7173) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM1(7173))))  severity failure;
	assert RAM1(7174) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM1(7174))))  severity failure;
	assert RAM1(7175) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM1(7175))))  severity failure;
	assert RAM1(7176) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM1(7176))))  severity failure;
	assert RAM1(7177) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM1(7177))))  severity failure;
	assert RAM1(7178) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM1(7178))))  severity failure;
	assert RAM1(7179) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM1(7179))))  severity failure;
	assert RAM1(7180) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM1(7180))))  severity failure;
	assert RAM1(7181) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM1(7181))))  severity failure;
	assert RAM1(7182) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM1(7182))))  severity failure;
	assert RAM1(7183) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM1(7183))))  severity failure;
	assert RAM1(7184) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM1(7184))))  severity failure;
	assert RAM1(7185) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM1(7185))))  severity failure;
	assert RAM1(7186) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM1(7186))))  severity failure;
	assert RAM1(7187) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM1(7187))))  severity failure;
	assert RAM1(7188) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM1(7188))))  severity failure;
	assert RAM1(7189) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM1(7189))))  severity failure;
	assert RAM1(7190) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM1(7190))))  severity failure;
	assert RAM1(7191) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM1(7191))))  severity failure;
	assert RAM1(7192) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM1(7192))))  severity failure;
	assert RAM1(7193) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM1(7193))))  severity failure;
	assert RAM1(7194) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM1(7194))))  severity failure;
	assert RAM1(7195) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM1(7195))))  severity failure;
	assert RAM1(7196) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM1(7196))))  severity failure;
	assert RAM1(7197) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM1(7197))))  severity failure;
	assert RAM1(7198) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM1(7198))))  severity failure;
	assert RAM1(7199) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM1(7199))))  severity failure;
	assert RAM1(7200) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM1(7200))))  severity failure;
	assert RAM1(7201) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM1(7201))))  severity failure;
	assert RAM1(7202) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM1(7202))))  severity failure;
	assert RAM1(7203) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM1(7203))))  severity failure;
	assert RAM1(7204) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM1(7204))))  severity failure;
	assert RAM1(7205) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM1(7205))))  severity failure;
	assert RAM1(7206) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM1(7206))))  severity failure;
	assert RAM1(7207) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM1(7207))))  severity failure;
	assert RAM1(7208) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM1(7208))))  severity failure;
	assert RAM1(7209) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM1(7209))))  severity failure;
	assert RAM1(7210) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM1(7210))))  severity failure;
	assert RAM1(7211) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM1(7211))))  severity failure;
	assert RAM1(7212) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM1(7212))))  severity failure;
	assert RAM1(7213) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM1(7213))))  severity failure;
	assert RAM1(7214) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM1(7214))))  severity failure;
	assert RAM1(7215) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM1(7215))))  severity failure;
	assert RAM1(7216) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM1(7216))))  severity failure;
	assert RAM1(7217) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM1(7217))))  severity failure;
	assert RAM1(7218) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM1(7218))))  severity failure;
	assert RAM1(7219) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM1(7219))))  severity failure;
	assert RAM1(7220) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM1(7220))))  severity failure;
	assert RAM1(7221) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM1(7221))))  severity failure;

	assert RAM2(1658) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM2(1658))))  severity failure;
	assert RAM2(1659) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM2(1659))))  severity failure;
	assert RAM2(1660) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM2(1660))))  severity failure;
	assert RAM2(1661) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM2(1661))))  severity failure;
	assert RAM2(1662) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM2(1662))))  severity failure;
	assert RAM2(1663) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM2(1663))))  severity failure;
	assert RAM2(1664) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM2(1664))))  severity failure;
	assert RAM2(1665) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM2(1665))))  severity failure;
	assert RAM2(1666) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM2(1666))))  severity failure;
	assert RAM2(1667) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM2(1667))))  severity failure;
	assert RAM2(1668) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM2(1668))))  severity failure;
	assert RAM2(1669) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM2(1669))))  severity failure;
	assert RAM2(1670) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM2(1670))))  severity failure;
	assert RAM2(1671) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM2(1671))))  severity failure;
	assert RAM2(1672) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM2(1672))))  severity failure;
	assert RAM2(1673) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM2(1673))))  severity failure;
	assert RAM2(1674) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM2(1674))))  severity failure;
	assert RAM2(1675) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM2(1675))))  severity failure;
	assert RAM2(1676) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM2(1676))))  severity failure;
	assert RAM2(1677) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM2(1677))))  severity failure;
	assert RAM2(1678) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM2(1678))))  severity failure;
	assert RAM2(1679) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM2(1679))))  severity failure;
	assert RAM2(1680) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM2(1680))))  severity failure;
	assert RAM2(1681) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM2(1681))))  severity failure;
	assert RAM2(1682) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM2(1682))))  severity failure;
	assert RAM2(1683) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM2(1683))))  severity failure;
	assert RAM2(1684) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM2(1684))))  severity failure;
	assert RAM2(1685) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM2(1685))))  severity failure;
	assert RAM2(1686) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM2(1686))))  severity failure;
	assert RAM2(1687) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM2(1687))))  severity failure;
	assert RAM2(1688) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM2(1688))))  severity failure;
	assert RAM2(1689) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM2(1689))))  severity failure;
	assert RAM2(1690) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM2(1690))))  severity failure;
	assert RAM2(1691) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM2(1691))))  severity failure;
	assert RAM2(1692) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM2(1692))))  severity failure;
	assert RAM2(1693) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM2(1693))))  severity failure;
	assert RAM2(1694) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM2(1694))))  severity failure;
	assert RAM2(1695) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM2(1695))))  severity failure;
	assert RAM2(1696) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM2(1696))))  severity failure;
	assert RAM2(1697) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM2(1697))))  severity failure;
	assert RAM2(1698) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM2(1698))))  severity failure;
	assert RAM2(1699) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM2(1699))))  severity failure;
	assert RAM2(1700) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM2(1700))))  severity failure;
	assert RAM2(1701) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM2(1701))))  severity failure;
	assert RAM2(1702) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM2(1702))))  severity failure;
	assert RAM2(1703) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM2(1703))))  severity failure;
	assert RAM2(1704) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM2(1704))))  severity failure;
	assert RAM2(1705) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM2(1705))))  severity failure;
	assert RAM2(1706) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM2(1706))))  severity failure;
	assert RAM2(1707) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM2(1707))))  severity failure;
	assert RAM2(1708) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM2(1708))))  severity failure;
	assert RAM2(1709) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM2(1709))))  severity failure;
	assert RAM2(1710) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM2(1710))))  severity failure;
	assert RAM2(1711) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM2(1711))))  severity failure;
	assert RAM2(1712) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM2(1712))))  severity failure;
	assert RAM2(1713) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM2(1713))))  severity failure;
	assert RAM2(1714) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM2(1714))))  severity failure;
	assert RAM2(1715) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM2(1715))))  severity failure;
	assert RAM2(1716) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM2(1716))))  severity failure;
	assert RAM2(1717) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM2(1717))))  severity failure;
	assert RAM2(1718) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM2(1718))))  severity failure;
	assert RAM2(1719) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM2(1719))))  severity failure;
	assert RAM2(1720) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM2(1720))))  severity failure;
	assert RAM2(1721) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM2(1721))))  severity failure;
	assert RAM2(1722) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM2(1722))))  severity failure;
	assert RAM2(1723) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM2(1723))))  severity failure;
	assert RAM2(1724) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM2(1724))))  severity failure;
	assert RAM2(1725) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM2(1725))))  severity failure;
	assert RAM2(1726) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM2(1726))))  severity failure;
	assert RAM2(1727) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM2(1727))))  severity failure;
	assert RAM2(1728) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM2(1728))))  severity failure;
	assert RAM2(1729) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM2(1729))))  severity failure;
	assert RAM2(1730) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM2(1730))))  severity failure;
	assert RAM2(1731) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM2(1731))))  severity failure;
	assert RAM2(1732) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM2(1732))))  severity failure;
	assert RAM2(1733) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM2(1733))))  severity failure;
	assert RAM2(1734) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM2(1734))))  severity failure;
	assert RAM2(1735) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM2(1735))))  severity failure;
	assert RAM2(1736) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM2(1736))))  severity failure;
	assert RAM2(1737) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM2(1737))))  severity failure;
	assert RAM2(1738) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM2(1738))))  severity failure;
	assert RAM2(1739) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM2(1739))))  severity failure;
	assert RAM2(1740) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM2(1740))))  severity failure;
	assert RAM2(1741) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM2(1741))))  severity failure;
	assert RAM2(1742) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM2(1742))))  severity failure;
	assert RAM2(1743) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM2(1743))))  severity failure;
	assert RAM2(1744) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM2(1744))))  severity failure;
	assert RAM2(1745) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM2(1745))))  severity failure;
	assert RAM2(1746) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM2(1746))))  severity failure;
	assert RAM2(1747) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM2(1747))))  severity failure;
	assert RAM2(1748) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM2(1748))))  severity failure;
	assert RAM2(1749) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM2(1749))))  severity failure;
	assert RAM2(1750) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM2(1750))))  severity failure;
	assert RAM2(1751) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM2(1751))))  severity failure;
	assert RAM2(1752) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM2(1752))))  severity failure;
	assert RAM2(1753) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM2(1753))))  severity failure;
	assert RAM2(1754) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM2(1754))))  severity failure;
	assert RAM2(1755) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM2(1755))))  severity failure;
	assert RAM2(1756) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM2(1756))))  severity failure;
	assert RAM2(1757) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM2(1757))))  severity failure;
	assert RAM2(1758) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM2(1758))))  severity failure;
	assert RAM2(1759) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM2(1759))))  severity failure;
	assert RAM2(1760) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM2(1760))))  severity failure;
	assert RAM2(1761) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM2(1761))))  severity failure;
	assert RAM2(1762) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM2(1762))))  severity failure;
	assert RAM2(1763) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM2(1763))))  severity failure;
	assert RAM2(1764) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM2(1764))))  severity failure;
	assert RAM2(1765) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM2(1765))))  severity failure;
	assert RAM2(1766) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM2(1766))))  severity failure;
	assert RAM2(1767) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM2(1767))))  severity failure;
	assert RAM2(1768) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM2(1768))))  severity failure;
	assert RAM2(1769) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM2(1769))))  severity failure;
	assert RAM2(1770) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM2(1770))))  severity failure;
	assert RAM2(1771) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM2(1771))))  severity failure;
	assert RAM2(1772) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM2(1772))))  severity failure;
	assert RAM2(1773) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM2(1773))))  severity failure;
	assert RAM2(1774) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM2(1774))))  severity failure;
	assert RAM2(1775) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM2(1775))))  severity failure;
	assert RAM2(1776) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM2(1776))))  severity failure;
	assert RAM2(1777) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM2(1777))))  severity failure;
	assert RAM2(1778) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM2(1778))))  severity failure;
	assert RAM2(1779) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM2(1779))))  severity failure;
	assert RAM2(1780) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM2(1780))))  severity failure;
	assert RAM2(1781) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM2(1781))))  severity failure;
	assert RAM2(1782) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM2(1782))))  severity failure;
	assert RAM2(1783) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM2(1783))))  severity failure;
	assert RAM2(1784) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM2(1784))))  severity failure;
	assert RAM2(1785) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM2(1785))))  severity failure;
	assert RAM2(1786) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM2(1786))))  severity failure;
	assert RAM2(1787) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM2(1787))))  severity failure;
	assert RAM2(1788) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM2(1788))))  severity failure;
	assert RAM2(1789) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM2(1789))))  severity failure;
	assert RAM2(1790) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM2(1790))))  severity failure;
	assert RAM2(1791) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM2(1791))))  severity failure;
	assert RAM2(1792) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM2(1792))))  severity failure;
	assert RAM2(1793) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM2(1793))))  severity failure;
	assert RAM2(1794) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM2(1794))))  severity failure;
	assert RAM2(1795) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM2(1795))))  severity failure;
	assert RAM2(1796) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM2(1796))))  severity failure;
	assert RAM2(1797) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM2(1797))))  severity failure;
	assert RAM2(1798) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM2(1798))))  severity failure;
	assert RAM2(1799) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM2(1799))))  severity failure;
	assert RAM2(1800) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM2(1800))))  severity failure;
	assert RAM2(1801) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM2(1801))))  severity failure;
	assert RAM2(1802) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM2(1802))))  severity failure;
	assert RAM2(1803) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM2(1803))))  severity failure;
	assert RAM2(1804) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM2(1804))))  severity failure;
	assert RAM2(1805) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM2(1805))))  severity failure;
	assert RAM2(1806) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM2(1806))))  severity failure;
	assert RAM2(1807) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM2(1807))))  severity failure;
	assert RAM2(1808) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM2(1808))))  severity failure;
	assert RAM2(1809) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM2(1809))))  severity failure;
	assert RAM2(1810) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM2(1810))))  severity failure;
	assert RAM2(1811) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM2(1811))))  severity failure;
	assert RAM2(1812) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM2(1812))))  severity failure;
	assert RAM2(1813) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM2(1813))))  severity failure;
	assert RAM2(1814) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM2(1814))))  severity failure;
	assert RAM2(1815) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM2(1815))))  severity failure;
	assert RAM2(1816) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM2(1816))))  severity failure;
	assert RAM2(1817) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM2(1817))))  severity failure;
	assert RAM2(1818) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM2(1818))))  severity failure;
	assert RAM2(1819) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM2(1819))))  severity failure;
	assert RAM2(1820) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM2(1820))))  severity failure;
	assert RAM2(1821) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM2(1821))))  severity failure;
	assert RAM2(1822) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM2(1822))))  severity failure;
	assert RAM2(1823) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM2(1823))))  severity failure;
	assert RAM2(1824) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM2(1824))))  severity failure;
	assert RAM2(1825) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM2(1825))))  severity failure;
	assert RAM2(1826) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM2(1826))))  severity failure;
	assert RAM2(1827) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM2(1827))))  severity failure;
	assert RAM2(1828) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM2(1828))))  severity failure;
	assert RAM2(1829) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM2(1829))))  severity failure;
	assert RAM2(1830) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM2(1830))))  severity failure;
	assert RAM2(1831) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM2(1831))))  severity failure;
	assert RAM2(1832) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM2(1832))))  severity failure;
	assert RAM2(1833) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM2(1833))))  severity failure;
	assert RAM2(1834) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM2(1834))))  severity failure;
	assert RAM2(1835) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM2(1835))))  severity failure;
	assert RAM2(1836) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM2(1836))))  severity failure;
	assert RAM2(1837) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM2(1837))))  severity failure;
	assert RAM2(1838) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM2(1838))))  severity failure;
	assert RAM2(1839) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM2(1839))))  severity failure;
	assert RAM2(1840) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM2(1840))))  severity failure;
	assert RAM2(1841) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM2(1841))))  severity failure;
	assert RAM2(1842) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM2(1842))))  severity failure;
	assert RAM2(1843) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM2(1843))))  severity failure;
	assert RAM2(1844) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM2(1844))))  severity failure;
	assert RAM2(1845) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM2(1845))))  severity failure;
	assert RAM2(1846) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM2(1846))))  severity failure;
	assert RAM2(1847) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM2(1847))))  severity failure;
	assert RAM2(1848) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM2(1848))))  severity failure;
	assert RAM2(1849) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM2(1849))))  severity failure;
	assert RAM2(1850) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM2(1850))))  severity failure;
	assert RAM2(1851) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM2(1851))))  severity failure;
	assert RAM2(1852) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM2(1852))))  severity failure;
	assert RAM2(1853) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM2(1853))))  severity failure;
	assert RAM2(1854) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM2(1854))))  severity failure;
	assert RAM2(1855) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM2(1855))))  severity failure;
	assert RAM2(1856) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM2(1856))))  severity failure;
	assert RAM2(1857) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM2(1857))))  severity failure;
	assert RAM2(1858) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM2(1858))))  severity failure;
	assert RAM2(1859) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM2(1859))))  severity failure;
	assert RAM2(1860) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM2(1860))))  severity failure;
	assert RAM2(1861) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM2(1861))))  severity failure;
	assert RAM2(1862) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM2(1862))))  severity failure;
	assert RAM2(1863) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM2(1863))))  severity failure;
	assert RAM2(1864) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM2(1864))))  severity failure;
	assert RAM2(1865) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM2(1865))))  severity failure;
	assert RAM2(1866) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM2(1866))))  severity failure;
	assert RAM2(1867) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM2(1867))))  severity failure;
	assert RAM2(1868) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM2(1868))))  severity failure;
	assert RAM2(1869) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM2(1869))))  severity failure;
	assert RAM2(1870) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM2(1870))))  severity failure;
	assert RAM2(1871) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM2(1871))))  severity failure;
	assert RAM2(1872) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM2(1872))))  severity failure;
	assert RAM2(1873) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM2(1873))))  severity failure;
	assert RAM2(1874) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM2(1874))))  severity failure;
	assert RAM2(1875) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM2(1875))))  severity failure;
	assert RAM2(1876) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM2(1876))))  severity failure;
	assert RAM2(1877) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM2(1877))))  severity failure;
	assert RAM2(1878) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM2(1878))))  severity failure;
	assert RAM2(1879) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM2(1879))))  severity failure;
	assert RAM2(1880) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM2(1880))))  severity failure;
	assert RAM2(1881) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM2(1881))))  severity failure;
	assert RAM2(1882) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM2(1882))))  severity failure;
	assert RAM2(1883) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM2(1883))))  severity failure;
	assert RAM2(1884) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM2(1884))))  severity failure;
	assert RAM2(1885) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM2(1885))))  severity failure;
	assert RAM2(1886) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM2(1886))))  severity failure;
	assert RAM2(1887) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM2(1887))))  severity failure;
	assert RAM2(1888) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM2(1888))))  severity failure;
	assert RAM2(1889) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM2(1889))))  severity failure;
	assert RAM2(1890) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM2(1890))))  severity failure;
	assert RAM2(1891) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM2(1891))))  severity failure;
	assert RAM2(1892) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM2(1892))))  severity failure;
	assert RAM2(1893) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM2(1893))))  severity failure;
	assert RAM2(1894) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM2(1894))))  severity failure;
	assert RAM2(1895) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM2(1895))))  severity failure;
	assert RAM2(1896) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM2(1896))))  severity failure;
	assert RAM2(1897) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM2(1897))))  severity failure;
	assert RAM2(1898) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM2(1898))))  severity failure;
	assert RAM2(1899) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM2(1899))))  severity failure;
	assert RAM2(1900) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM2(1900))))  severity failure;
	assert RAM2(1901) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM2(1901))))  severity failure;
	assert RAM2(1902) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM2(1902))))  severity failure;
	assert RAM2(1903) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM2(1903))))  severity failure;
	assert RAM2(1904) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM2(1904))))  severity failure;
	assert RAM2(1905) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM2(1905))))  severity failure;
	assert RAM2(1906) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM2(1906))))  severity failure;
	assert RAM2(1907) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM2(1907))))  severity failure;
	assert RAM2(1908) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM2(1908))))  severity failure;
	assert RAM2(1909) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM2(1909))))  severity failure;
	assert RAM2(1910) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM2(1910))))  severity failure;
	assert RAM2(1911) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM2(1911))))  severity failure;
	assert RAM2(1912) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM2(1912))))  severity failure;
	assert RAM2(1913) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM2(1913))))  severity failure;
	assert RAM2(1914) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM2(1914))))  severity failure;
	assert RAM2(1915) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM2(1915))))  severity failure;
	assert RAM2(1916) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM2(1916))))  severity failure;
	assert RAM2(1917) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM2(1917))))  severity failure;
	assert RAM2(1918) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM2(1918))))  severity failure;
	assert RAM2(1919) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM2(1919))))  severity failure;
	assert RAM2(1920) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM2(1920))))  severity failure;
	assert RAM2(1921) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM2(1921))))  severity failure;
	assert RAM2(1922) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM2(1922))))  severity failure;
	assert RAM2(1923) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM2(1923))))  severity failure;
	assert RAM2(1924) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM2(1924))))  severity failure;
	assert RAM2(1925) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM2(1925))))  severity failure;
	assert RAM2(1926) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM2(1926))))  severity failure;
	assert RAM2(1927) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM2(1927))))  severity failure;
	assert RAM2(1928) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM2(1928))))  severity failure;
	assert RAM2(1929) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM2(1929))))  severity failure;
	assert RAM2(1930) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM2(1930))))  severity failure;
	assert RAM2(1931) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM2(1931))))  severity failure;
	assert RAM2(1932) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM2(1932))))  severity failure;
	assert RAM2(1933) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM2(1933))))  severity failure;
	assert RAM2(1934) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM2(1934))))  severity failure;
	assert RAM2(1935) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM2(1935))))  severity failure;
	assert RAM2(1936) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM2(1936))))  severity failure;
	assert RAM2(1937) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM2(1937))))  severity failure;
	assert RAM2(1938) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM2(1938))))  severity failure;
	assert RAM2(1939) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM2(1939))))  severity failure;
	assert RAM2(1940) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM2(1940))))  severity failure;
	assert RAM2(1941) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM2(1941))))  severity failure;
	assert RAM2(1942) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM2(1942))))  severity failure;
	assert RAM2(1943) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM2(1943))))  severity failure;
	assert RAM2(1944) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM2(1944))))  severity failure;
	assert RAM2(1945) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM2(1945))))  severity failure;
	assert RAM2(1946) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM2(1946))))  severity failure;
	assert RAM2(1947) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM2(1947))))  severity failure;
	assert RAM2(1948) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM2(1948))))  severity failure;
	assert RAM2(1949) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM2(1949))))  severity failure;
	assert RAM2(1950) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM2(1950))))  severity failure;
	assert RAM2(1951) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM2(1951))))  severity failure;
	assert RAM2(1952) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM2(1952))))  severity failure;
	assert RAM2(1953) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM2(1953))))  severity failure;
	assert RAM2(1954) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM2(1954))))  severity failure;
	assert RAM2(1955) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM2(1955))))  severity failure;
	assert RAM2(1956) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM2(1956))))  severity failure;
	assert RAM2(1957) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM2(1957))))  severity failure;
	assert RAM2(1958) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM2(1958))))  severity failure;
	assert RAM2(1959) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM2(1959))))  severity failure;
	assert RAM2(1960) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM2(1960))))  severity failure;
	assert RAM2(1961) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM2(1961))))  severity failure;
	assert RAM2(1962) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM2(1962))))  severity failure;
	assert RAM2(1963) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM2(1963))))  severity failure;
	assert RAM2(1964) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM2(1964))))  severity failure;
	assert RAM2(1965) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM2(1965))))  severity failure;
	assert RAM2(1966) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM2(1966))))  severity failure;
	assert RAM2(1967) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM2(1967))))  severity failure;
	assert RAM2(1968) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM2(1968))))  severity failure;
	assert RAM2(1969) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM2(1969))))  severity failure;
	assert RAM2(1970) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM2(1970))))  severity failure;
	assert RAM2(1971) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM2(1971))))  severity failure;
	assert RAM2(1972) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM2(1972))))  severity failure;
	assert RAM2(1973) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM2(1973))))  severity failure;
	assert RAM2(1974) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM2(1974))))  severity failure;
	assert RAM2(1975) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM2(1975))))  severity failure;
	assert RAM2(1976) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM2(1976))))  severity failure;
	assert RAM2(1977) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM2(1977))))  severity failure;
	assert RAM2(1978) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM2(1978))))  severity failure;
	assert RAM2(1979) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM2(1979))))  severity failure;
	assert RAM2(1980) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM2(1980))))  severity failure;
	assert RAM2(1981) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM2(1981))))  severity failure;
	assert RAM2(1982) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM2(1982))))  severity failure;
	assert RAM2(1983) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM2(1983))))  severity failure;
	assert RAM2(1984) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM2(1984))))  severity failure;
	assert RAM2(1985) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM2(1985))))  severity failure;
	assert RAM2(1986) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM2(1986))))  severity failure;
	assert RAM2(1987) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM2(1987))))  severity failure;
	assert RAM2(1988) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM2(1988))))  severity failure;
	assert RAM2(1989) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM2(1989))))  severity failure;
	assert RAM2(1990) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM2(1990))))  severity failure;
	assert RAM2(1991) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM2(1991))))  severity failure;
	assert RAM2(1992) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM2(1992))))  severity failure;
	assert RAM2(1993) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM2(1993))))  severity failure;
	assert RAM2(1994) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM2(1994))))  severity failure;
	assert RAM2(1995) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM2(1995))))  severity failure;
	assert RAM2(1996) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM2(1996))))  severity failure;
	assert RAM2(1997) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM2(1997))))  severity failure;
	assert RAM2(1998) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM2(1998))))  severity failure;
	assert RAM2(1999) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM2(1999))))  severity failure;
	assert RAM2(2000) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM2(2000))))  severity failure;
	assert RAM2(2001) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM2(2001))))  severity failure;
	assert RAM2(2002) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM2(2002))))  severity failure;
	assert RAM2(2003) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM2(2003))))  severity failure;
	assert RAM2(2004) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM2(2004))))  severity failure;
	assert RAM2(2005) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM2(2005))))  severity failure;
	assert RAM2(2006) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM2(2006))))  severity failure;
	assert RAM2(2007) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM2(2007))))  severity failure;
	assert RAM2(2008) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM2(2008))))  severity failure;
	assert RAM2(2009) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM2(2009))))  severity failure;
	assert RAM2(2010) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM2(2010))))  severity failure;
	assert RAM2(2011) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM2(2011))))  severity failure;
	assert RAM2(2012) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM2(2012))))  severity failure;
	assert RAM2(2013) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM2(2013))))  severity failure;
	assert RAM2(2014) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM2(2014))))  severity failure;
	assert RAM2(2015) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM2(2015))))  severity failure;
	assert RAM2(2016) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM2(2016))))  severity failure;
	assert RAM2(2017) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM2(2017))))  severity failure;
	assert RAM2(2018) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM2(2018))))  severity failure;
	assert RAM2(2019) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM2(2019))))  severity failure;
	assert RAM2(2020) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM2(2020))))  severity failure;
	assert RAM2(2021) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM2(2021))))  severity failure;
	assert RAM2(2022) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM2(2022))))  severity failure;
	assert RAM2(2023) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM2(2023))))  severity failure;
	assert RAM2(2024) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM2(2024))))  severity failure;
	assert RAM2(2025) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM2(2025))))  severity failure;
	assert RAM2(2026) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM2(2026))))  severity failure;
	assert RAM2(2027) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM2(2027))))  severity failure;
	assert RAM2(2028) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM2(2028))))  severity failure;
	assert RAM2(2029) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM2(2029))))  severity failure;
	assert RAM2(2030) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM2(2030))))  severity failure;
	assert RAM2(2031) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM2(2031))))  severity failure;
	assert RAM2(2032) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM2(2032))))  severity failure;
	assert RAM2(2033) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM2(2033))))  severity failure;
	assert RAM2(2034) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM2(2034))))  severity failure;
	assert RAM2(2035) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM2(2035))))  severity failure;
	assert RAM2(2036) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM2(2036))))  severity failure;
	assert RAM2(2037) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM2(2037))))  severity failure;
	assert RAM2(2038) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM2(2038))))  severity failure;
	assert RAM2(2039) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM2(2039))))  severity failure;
	assert RAM2(2040) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM2(2040))))  severity failure;
	assert RAM2(2041) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM2(2041))))  severity failure;
	assert RAM2(2042) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM2(2042))))  severity failure;
	assert RAM2(2043) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM2(2043))))  severity failure;
	assert RAM2(2044) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM2(2044))))  severity failure;
	assert RAM2(2045) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM2(2045))))  severity failure;
	assert RAM2(2046) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM2(2046))))  severity failure;
	assert RAM2(2047) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM2(2047))))  severity failure;
	assert RAM2(2048) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM2(2048))))  severity failure;
	assert RAM2(2049) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM2(2049))))  severity failure;
	assert RAM2(2050) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM2(2050))))  severity failure;
	assert RAM2(2051) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM2(2051))))  severity failure;
	assert RAM2(2052) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM2(2052))))  severity failure;
	assert RAM2(2053) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM2(2053))))  severity failure;
	assert RAM2(2054) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM2(2054))))  severity failure;
	assert RAM2(2055) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM2(2055))))  severity failure;
	assert RAM2(2056) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM2(2056))))  severity failure;
	assert RAM2(2057) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM2(2057))))  severity failure;
	assert RAM2(2058) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM2(2058))))  severity failure;
	assert RAM2(2059) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM2(2059))))  severity failure;
	assert RAM2(2060) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM2(2060))))  severity failure;
	assert RAM2(2061) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM2(2061))))  severity failure;
	assert RAM2(2062) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM2(2062))))  severity failure;
	assert RAM2(2063) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM2(2063))))  severity failure;
	assert RAM2(2064) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM2(2064))))  severity failure;
	assert RAM2(2065) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM2(2065))))  severity failure;
	assert RAM2(2066) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM2(2066))))  severity failure;
	assert RAM2(2067) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM2(2067))))  severity failure;
	assert RAM2(2068) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM2(2068))))  severity failure;
	assert RAM2(2069) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM2(2069))))  severity failure;
	assert RAM2(2070) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM2(2070))))  severity failure;
	assert RAM2(2071) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM2(2071))))  severity failure;
	assert RAM2(2072) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM2(2072))))  severity failure;
	assert RAM2(2073) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM2(2073))))  severity failure;
	assert RAM2(2074) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM2(2074))))  severity failure;
	assert RAM2(2075) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM2(2075))))  severity failure;
	assert RAM2(2076) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM2(2076))))  severity failure;
	assert RAM2(2077) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM2(2077))))  severity failure;
	assert RAM2(2078) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM2(2078))))  severity failure;
	assert RAM2(2079) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM2(2079))))  severity failure;
	assert RAM2(2080) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM2(2080))))  severity failure;
	assert RAM2(2081) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM2(2081))))  severity failure;
	assert RAM2(2082) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM2(2082))))  severity failure;
	assert RAM2(2083) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM2(2083))))  severity failure;
	assert RAM2(2084) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM2(2084))))  severity failure;
	assert RAM2(2085) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM2(2085))))  severity failure;
	assert RAM2(2086) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM2(2086))))  severity failure;
	assert RAM2(2087) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM2(2087))))  severity failure;
	assert RAM2(2088) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM2(2088))))  severity failure;
	assert RAM2(2089) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM2(2089))))  severity failure;
	assert RAM2(2090) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM2(2090))))  severity failure;
	assert RAM2(2091) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM2(2091))))  severity failure;
	assert RAM2(2092) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM2(2092))))  severity failure;
	assert RAM2(2093) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM2(2093))))  severity failure;
	assert RAM2(2094) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM2(2094))))  severity failure;
	assert RAM2(2095) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM2(2095))))  severity failure;
	assert RAM2(2096) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM2(2096))))  severity failure;
	assert RAM2(2097) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM2(2097))))  severity failure;
	assert RAM2(2098) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM2(2098))))  severity failure;
	assert RAM2(2099) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM2(2099))))  severity failure;
	assert RAM2(2100) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM2(2100))))  severity failure;
	assert RAM2(2101) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM2(2101))))  severity failure;
	assert RAM2(2102) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM2(2102))))  severity failure;
	assert RAM2(2103) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM2(2103))))  severity failure;
	assert RAM2(2104) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM2(2104))))  severity failure;
	assert RAM2(2105) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM2(2105))))  severity failure;
	assert RAM2(2106) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM2(2106))))  severity failure;
	assert RAM2(2107) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM2(2107))))  severity failure;
	assert RAM2(2108) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM2(2108))))  severity failure;
	assert RAM2(2109) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM2(2109))))  severity failure;
	assert RAM2(2110) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM2(2110))))  severity failure;
	assert RAM2(2111) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM2(2111))))  severity failure;
	assert RAM2(2112) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM2(2112))))  severity failure;
	assert RAM2(2113) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM2(2113))))  severity failure;
	assert RAM2(2114) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM2(2114))))  severity failure;
	assert RAM2(2115) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM2(2115))))  severity failure;
	assert RAM2(2116) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM2(2116))))  severity failure;
	assert RAM2(2117) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM2(2117))))  severity failure;
	assert RAM2(2118) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM2(2118))))  severity failure;
	assert RAM2(2119) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM2(2119))))  severity failure;
	assert RAM2(2120) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM2(2120))))  severity failure;
	assert RAM2(2121) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM2(2121))))  severity failure;
	assert RAM2(2122) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM2(2122))))  severity failure;
	assert RAM2(2123) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM2(2123))))  severity failure;
	assert RAM2(2124) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM2(2124))))  severity failure;
	assert RAM2(2125) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM2(2125))))  severity failure;
	assert RAM2(2126) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM2(2126))))  severity failure;
	assert RAM2(2127) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM2(2127))))  severity failure;
	assert RAM2(2128) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM2(2128))))  severity failure;
	assert RAM2(2129) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM2(2129))))  severity failure;
	assert RAM2(2130) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM2(2130))))  severity failure;
	assert RAM2(2131) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM2(2131))))  severity failure;
	assert RAM2(2132) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM2(2132))))  severity failure;
	assert RAM2(2133) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM2(2133))))  severity failure;
	assert RAM2(2134) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM2(2134))))  severity failure;
	assert RAM2(2135) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM2(2135))))  severity failure;
	assert RAM2(2136) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM2(2136))))  severity failure;
	assert RAM2(2137) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM2(2137))))  severity failure;
	assert RAM2(2138) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM2(2138))))  severity failure;
	assert RAM2(2139) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM2(2139))))  severity failure;
	assert RAM2(2140) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM2(2140))))  severity failure;
	assert RAM2(2141) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM2(2141))))  severity failure;
	assert RAM2(2142) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM2(2142))))  severity failure;
	assert RAM2(2143) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM2(2143))))  severity failure;
	assert RAM2(2144) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM2(2144))))  severity failure;
	assert RAM2(2145) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM2(2145))))  severity failure;
	assert RAM2(2146) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM2(2146))))  severity failure;
	assert RAM2(2147) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM2(2147))))  severity failure;
	assert RAM2(2148) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM2(2148))))  severity failure;
	assert RAM2(2149) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM2(2149))))  severity failure;
	assert RAM2(2150) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM2(2150))))  severity failure;
	assert RAM2(2151) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM2(2151))))  severity failure;
	assert RAM2(2152) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM2(2152))))  severity failure;
	assert RAM2(2153) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM2(2153))))  severity failure;
	assert RAM2(2154) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM2(2154))))  severity failure;
	assert RAM2(2155) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM2(2155))))  severity failure;
	assert RAM2(2156) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM2(2156))))  severity failure;
	assert RAM2(2157) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM2(2157))))  severity failure;
	assert RAM2(2158) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM2(2158))))  severity failure;
	assert RAM2(2159) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM2(2159))))  severity failure;
	assert RAM2(2160) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM2(2160))))  severity failure;
	assert RAM2(2161) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM2(2161))))  severity failure;
	assert RAM2(2162) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM2(2162))))  severity failure;
	assert RAM2(2163) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM2(2163))))  severity failure;
	assert RAM2(2164) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM2(2164))))  severity failure;
	assert RAM2(2165) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM2(2165))))  severity failure;
	assert RAM2(2166) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM2(2166))))  severity failure;
	assert RAM2(2167) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM2(2167))))  severity failure;
	assert RAM2(2168) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM2(2168))))  severity failure;
	assert RAM2(2169) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM2(2169))))  severity failure;
	assert RAM2(2170) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM2(2170))))  severity failure;
	assert RAM2(2171) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM2(2171))))  severity failure;
	assert RAM2(2172) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM2(2172))))  severity failure;
	assert RAM2(2173) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM2(2173))))  severity failure;
	assert RAM2(2174) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM2(2174))))  severity failure;
	assert RAM2(2175) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM2(2175))))  severity failure;
	assert RAM2(2176) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM2(2176))))  severity failure;
	assert RAM2(2177) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM2(2177))))  severity failure;
	assert RAM2(2178) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM2(2178))))  severity failure;
	assert RAM2(2179) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM2(2179))))  severity failure;
	assert RAM2(2180) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM2(2180))))  severity failure;
	assert RAM2(2181) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM2(2181))))  severity failure;
	assert RAM2(2182) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM2(2182))))  severity failure;
	assert RAM2(2183) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM2(2183))))  severity failure;
	assert RAM2(2184) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM2(2184))))  severity failure;
	assert RAM2(2185) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM2(2185))))  severity failure;
	assert RAM2(2186) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM2(2186))))  severity failure;
	assert RAM2(2187) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM2(2187))))  severity failure;
	assert RAM2(2188) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM2(2188))))  severity failure;
	assert RAM2(2189) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM2(2189))))  severity failure;
	assert RAM2(2190) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM2(2190))))  severity failure;
	assert RAM2(2191) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM2(2191))))  severity failure;
	assert RAM2(2192) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM2(2192))))  severity failure;
	assert RAM2(2193) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM2(2193))))  severity failure;
	assert RAM2(2194) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM2(2194))))  severity failure;
	assert RAM2(2195) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM2(2195))))  severity failure;
	assert RAM2(2196) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM2(2196))))  severity failure;
	assert RAM2(2197) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM2(2197))))  severity failure;
	assert RAM2(2198) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM2(2198))))  severity failure;
	assert RAM2(2199) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM2(2199))))  severity failure;
	assert RAM2(2200) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM2(2200))))  severity failure;
	assert RAM2(2201) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM2(2201))))  severity failure;
	assert RAM2(2202) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM2(2202))))  severity failure;
	assert RAM2(2203) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM2(2203))))  severity failure;
	assert RAM2(2204) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM2(2204))))  severity failure;
	assert RAM2(2205) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM2(2205))))  severity failure;
	assert RAM2(2206) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM2(2206))))  severity failure;
	assert RAM2(2207) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM2(2207))))  severity failure;
	assert RAM2(2208) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM2(2208))))  severity failure;
	assert RAM2(2209) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM2(2209))))  severity failure;
	assert RAM2(2210) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM2(2210))))  severity failure;
	assert RAM2(2211) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM2(2211))))  severity failure;
	assert RAM2(2212) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM2(2212))))  severity failure;
	assert RAM2(2213) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM2(2213))))  severity failure;
	assert RAM2(2214) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM2(2214))))  severity failure;
	assert RAM2(2215) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM2(2215))))  severity failure;
	assert RAM2(2216) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM2(2216))))  severity failure;
	assert RAM2(2217) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM2(2217))))  severity failure;
	assert RAM2(2218) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM2(2218))))  severity failure;
	assert RAM2(2219) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM2(2219))))  severity failure;
	assert RAM2(2220) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM2(2220))))  severity failure;
	assert RAM2(2221) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM2(2221))))  severity failure;
	assert RAM2(2222) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM2(2222))))  severity failure;
	assert RAM2(2223) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM2(2223))))  severity failure;
	assert RAM2(2224) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM2(2224))))  severity failure;
	assert RAM2(2225) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM2(2225))))  severity failure;
	assert RAM2(2226) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM2(2226))))  severity failure;
	assert RAM2(2227) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM2(2227))))  severity failure;
	assert RAM2(2228) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM2(2228))))  severity failure;
	assert RAM2(2229) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM2(2229))))  severity failure;
	assert RAM2(2230) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM2(2230))))  severity failure;
	assert RAM2(2231) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM2(2231))))  severity failure;
	assert RAM2(2232) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM2(2232))))  severity failure;
	assert RAM2(2233) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM2(2233))))  severity failure;
	assert RAM2(2234) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM2(2234))))  severity failure;
	assert RAM2(2235) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM2(2235))))  severity failure;
	assert RAM2(2236) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM2(2236))))  severity failure;
	assert RAM2(2237) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM2(2237))))  severity failure;
	assert RAM2(2238) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM2(2238))))  severity failure;
	assert RAM2(2239) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM2(2239))))  severity failure;
	assert RAM2(2240) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM2(2240))))  severity failure;
	assert RAM2(2241) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM2(2241))))  severity failure;
	assert RAM2(2242) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM2(2242))))  severity failure;
	assert RAM2(2243) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM2(2243))))  severity failure;
	assert RAM2(2244) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM2(2244))))  severity failure;
	assert RAM2(2245) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM2(2245))))  severity failure;
	assert RAM2(2246) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM2(2246))))  severity failure;
	assert RAM2(2247) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM2(2247))))  severity failure;
	assert RAM2(2248) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM2(2248))))  severity failure;
	assert RAM2(2249) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM2(2249))))  severity failure;
	assert RAM2(2250) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM2(2250))))  severity failure;
	assert RAM2(2251) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM2(2251))))  severity failure;
	assert RAM2(2252) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM2(2252))))  severity failure;
	assert RAM2(2253) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM2(2253))))  severity failure;
	assert RAM2(2254) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM2(2254))))  severity failure;
	assert RAM2(2255) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM2(2255))))  severity failure;
	assert RAM2(2256) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM2(2256))))  severity failure;
	assert RAM2(2257) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM2(2257))))  severity failure;
	assert RAM2(2258) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM2(2258))))  severity failure;
	assert RAM2(2259) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM2(2259))))  severity failure;
	assert RAM2(2260) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM2(2260))))  severity failure;
	assert RAM2(2261) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM2(2261))))  severity failure;
	assert RAM2(2262) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM2(2262))))  severity failure;
	assert RAM2(2263) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM2(2263))))  severity failure;
	assert RAM2(2264) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM2(2264))))  severity failure;
	assert RAM2(2265) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM2(2265))))  severity failure;
	assert RAM2(2266) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM2(2266))))  severity failure;
	assert RAM2(2267) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM2(2267))))  severity failure;
	assert RAM2(2268) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM2(2268))))  severity failure;
	assert RAM2(2269) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM2(2269))))  severity failure;
	assert RAM2(2270) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM2(2270))))  severity failure;
	assert RAM2(2271) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM2(2271))))  severity failure;
	assert RAM2(2272) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM2(2272))))  severity failure;
	assert RAM2(2273) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM2(2273))))  severity failure;
	assert RAM2(2274) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM2(2274))))  severity failure;
	assert RAM2(2275) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM2(2275))))  severity failure;
	assert RAM2(2276) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM2(2276))))  severity failure;
	assert RAM2(2277) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM2(2277))))  severity failure;
	assert RAM2(2278) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM2(2278))))  severity failure;
	assert RAM2(2279) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM2(2279))))  severity failure;
	assert RAM2(2280) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM2(2280))))  severity failure;
	assert RAM2(2281) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM2(2281))))  severity failure;
	assert RAM2(2282) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM2(2282))))  severity failure;
	assert RAM2(2283) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM2(2283))))  severity failure;
	assert RAM2(2284) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM2(2284))))  severity failure;
	assert RAM2(2285) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM2(2285))))  severity failure;
	assert RAM2(2286) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM2(2286))))  severity failure;
	assert RAM2(2287) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM2(2287))))  severity failure;
	assert RAM2(2288) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM2(2288))))  severity failure;
	assert RAM2(2289) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM2(2289))))  severity failure;
	assert RAM2(2290) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM2(2290))))  severity failure;
	assert RAM2(2291) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM2(2291))))  severity failure;
	assert RAM2(2292) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM2(2292))))  severity failure;
	assert RAM2(2293) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM2(2293))))  severity failure;
	assert RAM2(2294) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM2(2294))))  severity failure;
	assert RAM2(2295) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM2(2295))))  severity failure;
	assert RAM2(2296) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM2(2296))))  severity failure;
	assert RAM2(2297) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM2(2297))))  severity failure;
	assert RAM2(2298) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM2(2298))))  severity failure;
	assert RAM2(2299) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM2(2299))))  severity failure;
	assert RAM2(2300) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM2(2300))))  severity failure;
	assert RAM2(2301) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM2(2301))))  severity failure;
	assert RAM2(2302) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM2(2302))))  severity failure;
	assert RAM2(2303) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM2(2303))))  severity failure;
	assert RAM2(2304) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM2(2304))))  severity failure;
	assert RAM2(2305) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM2(2305))))  severity failure;
	assert RAM2(2306) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM2(2306))))  severity failure;
	assert RAM2(2307) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM2(2307))))  severity failure;
	assert RAM2(2308) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM2(2308))))  severity failure;
	assert RAM2(2309) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM2(2309))))  severity failure;
	assert RAM2(2310) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM2(2310))))  severity failure;
	assert RAM2(2311) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM2(2311))))  severity failure;
	assert RAM2(2312) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM2(2312))))  severity failure;
	assert RAM2(2313) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM2(2313))))  severity failure;
	assert RAM2(2314) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM2(2314))))  severity failure;
	assert RAM2(2315) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM2(2315))))  severity failure;
	assert RAM2(2316) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM2(2316))))  severity failure;
	assert RAM2(2317) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM2(2317))))  severity failure;
	assert RAM2(2318) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM2(2318))))  severity failure;
	assert RAM2(2319) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM2(2319))))  severity failure;
	assert RAM2(2320) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM2(2320))))  severity failure;
	assert RAM2(2321) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM2(2321))))  severity failure;
	assert RAM2(2322) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM2(2322))))  severity failure;
	assert RAM2(2323) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM2(2323))))  severity failure;
	assert RAM2(2324) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM2(2324))))  severity failure;
	assert RAM2(2325) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM2(2325))))  severity failure;
	assert RAM2(2326) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM2(2326))))  severity failure;
	assert RAM2(2327) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM2(2327))))  severity failure;
	assert RAM2(2328) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM2(2328))))  severity failure;
	assert RAM2(2329) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM2(2329))))  severity failure;
	assert RAM2(2330) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM2(2330))))  severity failure;
	assert RAM2(2331) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM2(2331))))  severity failure;
	assert RAM2(2332) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM2(2332))))  severity failure;
	assert RAM2(2333) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM2(2333))))  severity failure;
	assert RAM2(2334) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM2(2334))))  severity failure;
	assert RAM2(2335) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM2(2335))))  severity failure;
	assert RAM2(2336) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM2(2336))))  severity failure;
	assert RAM2(2337) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM2(2337))))  severity failure;
	assert RAM2(2338) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM2(2338))))  severity failure;
	assert RAM2(2339) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM2(2339))))  severity failure;
	assert RAM2(2340) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM2(2340))))  severity failure;
	assert RAM2(2341) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM2(2341))))  severity failure;
	assert RAM2(2342) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM2(2342))))  severity failure;
	assert RAM2(2343) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM2(2343))))  severity failure;
	assert RAM2(2344) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM2(2344))))  severity failure;
	assert RAM2(2345) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM2(2345))))  severity failure;
	assert RAM2(2346) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM2(2346))))  severity failure;
	assert RAM2(2347) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM2(2347))))  severity failure;
	assert RAM2(2348) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM2(2348))))  severity failure;
	assert RAM2(2349) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM2(2349))))  severity failure;
	assert RAM2(2350) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM2(2350))))  severity failure;
	assert RAM2(2351) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM2(2351))))  severity failure;
	assert RAM2(2352) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM2(2352))))  severity failure;
	assert RAM2(2353) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM2(2353))))  severity failure;
	assert RAM2(2354) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM2(2354))))  severity failure;
	assert RAM2(2355) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM2(2355))))  severity failure;
	assert RAM2(2356) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM2(2356))))  severity failure;
	assert RAM2(2357) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM2(2357))))  severity failure;
	assert RAM2(2358) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM2(2358))))  severity failure;
	assert RAM2(2359) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM2(2359))))  severity failure;
	assert RAM2(2360) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM2(2360))))  severity failure;
	assert RAM2(2361) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM2(2361))))  severity failure;
	assert RAM2(2362) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM2(2362))))  severity failure;
	assert RAM2(2363) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM2(2363))))  severity failure;
	assert RAM2(2364) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM2(2364))))  severity failure;
	assert RAM2(2365) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM2(2365))))  severity failure;
	assert RAM2(2366) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM2(2366))))  severity failure;
	assert RAM2(2367) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM2(2367))))  severity failure;
	assert RAM2(2368) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM2(2368))))  severity failure;
	assert RAM2(2369) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM2(2369))))  severity failure;
	assert RAM2(2370) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM2(2370))))  severity failure;
	assert RAM2(2371) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM2(2371))))  severity failure;
	assert RAM2(2372) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM2(2372))))  severity failure;
	assert RAM2(2373) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM2(2373))))  severity failure;
	assert RAM2(2374) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM2(2374))))  severity failure;
	assert RAM2(2375) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM2(2375))))  severity failure;
	assert RAM2(2376) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM2(2376))))  severity failure;
	assert RAM2(2377) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM2(2377))))  severity failure;
	assert RAM2(2378) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM2(2378))))  severity failure;
	assert RAM2(2379) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM2(2379))))  severity failure;
	assert RAM2(2380) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM2(2380))))  severity failure;
	assert RAM2(2381) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM2(2381))))  severity failure;
	assert RAM2(2382) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM2(2382))))  severity failure;
	assert RAM2(2383) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM2(2383))))  severity failure;
	assert RAM2(2384) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM2(2384))))  severity failure;
	assert RAM2(2385) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM2(2385))))  severity failure;
	assert RAM2(2386) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM2(2386))))  severity failure;
	assert RAM2(2387) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM2(2387))))  severity failure;
	assert RAM2(2388) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM2(2388))))  severity failure;
	assert RAM2(2389) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM2(2389))))  severity failure;
	assert RAM2(2390) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM2(2390))))  severity failure;
	assert RAM2(2391) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM2(2391))))  severity failure;
	assert RAM2(2392) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM2(2392))))  severity failure;
	assert RAM2(2393) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM2(2393))))  severity failure;
	assert RAM2(2394) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM2(2394))))  severity failure;
	assert RAM2(2395) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM2(2395))))  severity failure;
	assert RAM2(2396) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM2(2396))))  severity failure;
	assert RAM2(2397) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM2(2397))))  severity failure;
	assert RAM2(2398) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM2(2398))))  severity failure;
	assert RAM2(2399) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM2(2399))))  severity failure;
	assert RAM2(2400) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM2(2400))))  severity failure;
	assert RAM2(2401) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM2(2401))))  severity failure;
	assert RAM2(2402) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM2(2402))))  severity failure;
	assert RAM2(2403) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM2(2403))))  severity failure;
	assert RAM2(2404) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM2(2404))))  severity failure;
	assert RAM2(2405) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM2(2405))))  severity failure;
	assert RAM2(2406) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM2(2406))))  severity failure;
	assert RAM2(2407) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM2(2407))))  severity failure;
	assert RAM2(2408) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM2(2408))))  severity failure;
	assert RAM2(2409) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM2(2409))))  severity failure;
	assert RAM2(2410) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM2(2410))))  severity failure;
	assert RAM2(2411) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM2(2411))))  severity failure;
	assert RAM2(2412) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM2(2412))))  severity failure;
	assert RAM2(2413) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM2(2413))))  severity failure;
	assert RAM2(2414) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM2(2414))))  severity failure;
	assert RAM2(2415) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM2(2415))))  severity failure;
	assert RAM2(2416) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM2(2416))))  severity failure;
	assert RAM2(2417) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM2(2417))))  severity failure;
	assert RAM2(2418) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM2(2418))))  severity failure;
	assert RAM2(2419) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM2(2419))))  severity failure;
	assert RAM2(2420) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM2(2420))))  severity failure;
	assert RAM2(2421) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM2(2421))))  severity failure;
	assert RAM2(2422) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM2(2422))))  severity failure;
	assert RAM2(2423) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM2(2423))))  severity failure;
	assert RAM2(2424) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM2(2424))))  severity failure;
	assert RAM2(2425) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM2(2425))))  severity failure;
	assert RAM2(2426) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM2(2426))))  severity failure;
	assert RAM2(2427) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM2(2427))))  severity failure;
	assert RAM2(2428) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM2(2428))))  severity failure;
	assert RAM2(2429) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM2(2429))))  severity failure;
	assert RAM2(2430) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM2(2430))))  severity failure;
	assert RAM2(2431) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM2(2431))))  severity failure;
	assert RAM2(2432) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM2(2432))))  severity failure;
	assert RAM2(2433) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM2(2433))))  severity failure;
	assert RAM2(2434) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM2(2434))))  severity failure;
	assert RAM2(2435) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM2(2435))))  severity failure;
	assert RAM2(2436) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM2(2436))))  severity failure;
	assert RAM2(2437) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM2(2437))))  severity failure;
	assert RAM2(2438) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM2(2438))))  severity failure;
	assert RAM2(2439) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM2(2439))))  severity failure;
	assert RAM2(2440) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM2(2440))))  severity failure;
	assert RAM2(2441) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM2(2441))))  severity failure;
	assert RAM2(2442) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM2(2442))))  severity failure;
	assert RAM2(2443) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM2(2443))))  severity failure;
	assert RAM2(2444) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM2(2444))))  severity failure;
	assert RAM2(2445) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM2(2445))))  severity failure;
	assert RAM2(2446) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM2(2446))))  severity failure;
	assert RAM2(2447) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM2(2447))))  severity failure;
	assert RAM2(2448) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM2(2448))))  severity failure;
	assert RAM2(2449) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM2(2449))))  severity failure;
	assert RAM2(2450) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM2(2450))))  severity failure;
	assert RAM2(2451) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM2(2451))))  severity failure;
	assert RAM2(2452) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM2(2452))))  severity failure;
	assert RAM2(2453) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM2(2453))))  severity failure;
	assert RAM2(2454) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM2(2454))))  severity failure;
	assert RAM2(2455) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM2(2455))))  severity failure;
	assert RAM2(2456) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM2(2456))))  severity failure;
	assert RAM2(2457) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM2(2457))))  severity failure;
	assert RAM2(2458) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM2(2458))))  severity failure;
	assert RAM2(2459) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM2(2459))))  severity failure;
	assert RAM2(2460) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM2(2460))))  severity failure;
	assert RAM2(2461) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM2(2461))))  severity failure;
	assert RAM2(2462) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM2(2462))))  severity failure;
	assert RAM2(2463) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM2(2463))))  severity failure;
	assert RAM2(2464) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM2(2464))))  severity failure;
	assert RAM2(2465) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM2(2465))))  severity failure;
	assert RAM2(2466) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM2(2466))))  severity failure;
	assert RAM2(2467) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM2(2467))))  severity failure;
	assert RAM2(2468) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM2(2468))))  severity failure;
	assert RAM2(2469) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM2(2469))))  severity failure;
	assert RAM2(2470) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM2(2470))))  severity failure;
	assert RAM2(2471) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM2(2471))))  severity failure;
	assert RAM2(2472) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM2(2472))))  severity failure;
	assert RAM2(2473) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM2(2473))))  severity failure;
	assert RAM2(2474) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM2(2474))))  severity failure;
	assert RAM2(2475) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM2(2475))))  severity failure;
	assert RAM2(2476) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM2(2476))))  severity failure;
	assert RAM2(2477) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM2(2477))))  severity failure;
	assert RAM2(2478) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM2(2478))))  severity failure;
	assert RAM2(2479) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM2(2479))))  severity failure;
	assert RAM2(2480) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM2(2480))))  severity failure;
	assert RAM2(2481) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM2(2481))))  severity failure;
	assert RAM2(2482) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM2(2482))))  severity failure;
	assert RAM2(2483) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM2(2483))))  severity failure;
	assert RAM2(2484) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM2(2484))))  severity failure;
	assert RAM2(2485) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM2(2485))))  severity failure;
	assert RAM2(2486) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM2(2486))))  severity failure;
	assert RAM2(2487) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM2(2487))))  severity failure;
	assert RAM2(2488) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM2(2488))))  severity failure;
	assert RAM2(2489) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM2(2489))))  severity failure;
	assert RAM2(2490) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM2(2490))))  severity failure;
	assert RAM2(2491) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM2(2491))))  severity failure;
	assert RAM2(2492) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM2(2492))))  severity failure;
	assert RAM2(2493) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM2(2493))))  severity failure;
	assert RAM2(2494) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM2(2494))))  severity failure;
	assert RAM2(2495) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM2(2495))))  severity failure;
	assert RAM2(2496) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM2(2496))))  severity failure;
	assert RAM2(2497) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM2(2497))))  severity failure;
	assert RAM2(2498) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM2(2498))))  severity failure;
	assert RAM2(2499) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM2(2499))))  severity failure;
	assert RAM2(2500) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM2(2500))))  severity failure;
	assert RAM2(2501) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM2(2501))))  severity failure;
	assert RAM2(2502) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM2(2502))))  severity failure;
	assert RAM2(2503) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM2(2503))))  severity failure;
	assert RAM2(2504) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM2(2504))))  severity failure;
	assert RAM2(2505) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM2(2505))))  severity failure;
	assert RAM2(2506) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM2(2506))))  severity failure;
	assert RAM2(2507) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM2(2507))))  severity failure;
	assert RAM2(2508) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM2(2508))))  severity failure;
	assert RAM2(2509) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM2(2509))))  severity failure;
	assert RAM2(2510) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM2(2510))))  severity failure;
	assert RAM2(2511) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM2(2511))))  severity failure;
	assert RAM2(2512) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM2(2512))))  severity failure;
	assert RAM2(2513) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM2(2513))))  severity failure;
	assert RAM2(2514) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM2(2514))))  severity failure;
	assert RAM2(2515) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM2(2515))))  severity failure;
	assert RAM2(2516) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM2(2516))))  severity failure;
	assert RAM2(2517) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM2(2517))))  severity failure;
	assert RAM2(2518) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM2(2518))))  severity failure;
	assert RAM2(2519) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM2(2519))))  severity failure;
	assert RAM2(2520) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM2(2520))))  severity failure;
	assert RAM2(2521) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM2(2521))))  severity failure;
	assert RAM2(2522) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM2(2522))))  severity failure;
	assert RAM2(2523) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM2(2523))))  severity failure;
	assert RAM2(2524) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM2(2524))))  severity failure;
	assert RAM2(2525) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM2(2525))))  severity failure;
	assert RAM2(2526) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM2(2526))))  severity failure;
	assert RAM2(2527) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM2(2527))))  severity failure;
	assert RAM2(2528) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM2(2528))))  severity failure;
	assert RAM2(2529) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM2(2529))))  severity failure;
	assert RAM2(2530) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM2(2530))))  severity failure;
	assert RAM2(2531) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM2(2531))))  severity failure;
	assert RAM2(2532) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM2(2532))))  severity failure;
	assert RAM2(2533) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM2(2533))))  severity failure;
	assert RAM2(2534) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM2(2534))))  severity failure;
	assert RAM2(2535) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM2(2535))))  severity failure;
	assert RAM2(2536) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM2(2536))))  severity failure;
	assert RAM2(2537) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM2(2537))))  severity failure;
	assert RAM2(2538) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM2(2538))))  severity failure;
	assert RAM2(2539) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM2(2539))))  severity failure;
	assert RAM2(2540) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM2(2540))))  severity failure;
	assert RAM2(2541) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM2(2541))))  severity failure;
	assert RAM2(2542) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM2(2542))))  severity failure;
	assert RAM2(2543) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM2(2543))))  severity failure;
	assert RAM2(2544) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM2(2544))))  severity failure;
	assert RAM2(2545) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM2(2545))))  severity failure;
	assert RAM2(2546) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM2(2546))))  severity failure;
	assert RAM2(2547) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM2(2547))))  severity failure;
	assert RAM2(2548) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM2(2548))))  severity failure;
	assert RAM2(2549) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM2(2549))))  severity failure;
	assert RAM2(2550) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM2(2550))))  severity failure;
	assert RAM2(2551) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM2(2551))))  severity failure;
	assert RAM2(2552) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM2(2552))))  severity failure;
	assert RAM2(2553) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM2(2553))))  severity failure;
	assert RAM2(2554) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM2(2554))))  severity failure;
	assert RAM2(2555) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM2(2555))))  severity failure;
	assert RAM2(2556) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM2(2556))))  severity failure;
	assert RAM2(2557) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM2(2557))))  severity failure;
	assert RAM2(2558) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM2(2558))))  severity failure;
	assert RAM2(2559) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM2(2559))))  severity failure;
	assert RAM2(2560) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM2(2560))))  severity failure;
	assert RAM2(2561) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM2(2561))))  severity failure;
	assert RAM2(2562) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM2(2562))))  severity failure;
	assert RAM2(2563) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM2(2563))))  severity failure;
	assert RAM2(2564) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM2(2564))))  severity failure;
	assert RAM2(2565) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM2(2565))))  severity failure;
	assert RAM2(2566) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM2(2566))))  severity failure;
	assert RAM2(2567) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM2(2567))))  severity failure;
	assert RAM2(2568) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM2(2568))))  severity failure;
	assert RAM2(2569) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM2(2569))))  severity failure;
	assert RAM2(2570) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM2(2570))))  severity failure;
	assert RAM2(2571) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM2(2571))))  severity failure;
	assert RAM2(2572) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM2(2572))))  severity failure;
	assert RAM2(2573) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM2(2573))))  severity failure;
	assert RAM2(2574) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM2(2574))))  severity failure;
	assert RAM2(2575) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM2(2575))))  severity failure;
	assert RAM2(2576) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM2(2576))))  severity failure;
	assert RAM2(2577) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM2(2577))))  severity failure;
	assert RAM2(2578) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM2(2578))))  severity failure;
	assert RAM2(2579) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM2(2579))))  severity failure;
	assert RAM2(2580) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM2(2580))))  severity failure;
	assert RAM2(2581) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM2(2581))))  severity failure;
	assert RAM2(2582) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM2(2582))))  severity failure;
	assert RAM2(2583) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM2(2583))))  severity failure;
	assert RAM2(2584) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM2(2584))))  severity failure;
	assert RAM2(2585) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM2(2585))))  severity failure;
	assert RAM2(2586) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM2(2586))))  severity failure;
	assert RAM2(2587) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM2(2587))))  severity failure;
	assert RAM2(2588) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM2(2588))))  severity failure;
	assert RAM2(2589) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM2(2589))))  severity failure;
	assert RAM2(2590) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM2(2590))))  severity failure;
	assert RAM2(2591) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM2(2591))))  severity failure;
	assert RAM2(2592) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM2(2592))))  severity failure;
	assert RAM2(2593) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM2(2593))))  severity failure;
	assert RAM2(2594) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM2(2594))))  severity failure;
	assert RAM2(2595) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM2(2595))))  severity failure;
	assert RAM2(2596) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM2(2596))))  severity failure;
	assert RAM2(2597) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM2(2597))))  severity failure;
	assert RAM2(2598) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM2(2598))))  severity failure;
	assert RAM2(2599) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM2(2599))))  severity failure;
	assert RAM2(2600) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM2(2600))))  severity failure;
	assert RAM2(2601) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM2(2601))))  severity failure;
	assert RAM2(2602) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM2(2602))))  severity failure;
	assert RAM2(2603) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM2(2603))))  severity failure;
	assert RAM2(2604) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM2(2604))))  severity failure;
	assert RAM2(2605) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM2(2605))))  severity failure;
	assert RAM2(2606) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM2(2606))))  severity failure;
	assert RAM2(2607) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM2(2607))))  severity failure;
	assert RAM2(2608) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM2(2608))))  severity failure;
	assert RAM2(2609) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM2(2609))))  severity failure;
	assert RAM2(2610) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM2(2610))))  severity failure;
	assert RAM2(2611) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM2(2611))))  severity failure;
	assert RAM2(2612) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM2(2612))))  severity failure;
	assert RAM2(2613) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM2(2613))))  severity failure;
	assert RAM2(2614) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM2(2614))))  severity failure;
	assert RAM2(2615) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM2(2615))))  severity failure;
	assert RAM2(2616) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM2(2616))))  severity failure;
	assert RAM2(2617) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM2(2617))))  severity failure;
	assert RAM2(2618) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM2(2618))))  severity failure;
	assert RAM2(2619) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM2(2619))))  severity failure;
	assert RAM2(2620) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM2(2620))))  severity failure;
	assert RAM2(2621) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM2(2621))))  severity failure;
	assert RAM2(2622) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM2(2622))))  severity failure;
	assert RAM2(2623) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM2(2623))))  severity failure;
	assert RAM2(2624) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM2(2624))))  severity failure;
	assert RAM2(2625) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM2(2625))))  severity failure;
	assert RAM2(2626) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM2(2626))))  severity failure;
	assert RAM2(2627) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM2(2627))))  severity failure;
	assert RAM2(2628) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM2(2628))))  severity failure;
	assert RAM2(2629) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM2(2629))))  severity failure;
	assert RAM2(2630) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM2(2630))))  severity failure;
	assert RAM2(2631) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM2(2631))))  severity failure;
	assert RAM2(2632) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM2(2632))))  severity failure;
	assert RAM2(2633) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM2(2633))))  severity failure;
	assert RAM2(2634) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM2(2634))))  severity failure;
	assert RAM2(2635) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM2(2635))))  severity failure;
	assert RAM2(2636) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM2(2636))))  severity failure;
	assert RAM2(2637) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM2(2637))))  severity failure;
	assert RAM2(2638) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM2(2638))))  severity failure;
	assert RAM2(2639) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM2(2639))))  severity failure;
	assert RAM2(2640) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM2(2640))))  severity failure;
	assert RAM2(2641) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM2(2641))))  severity failure;
	assert RAM2(2642) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM2(2642))))  severity failure;
	assert RAM2(2643) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM2(2643))))  severity failure;
	assert RAM2(2644) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM2(2644))))  severity failure;
	assert RAM2(2645) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM2(2645))))  severity failure;
	assert RAM2(2646) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM2(2646))))  severity failure;
	assert RAM2(2647) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM2(2647))))  severity failure;
	assert RAM2(2648) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM2(2648))))  severity failure;
	assert RAM2(2649) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM2(2649))))  severity failure;
	assert RAM2(2650) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM2(2650))))  severity failure;
	assert RAM2(2651) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM2(2651))))  severity failure;
	assert RAM2(2652) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM2(2652))))  severity failure;
	assert RAM2(2653) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM2(2653))))  severity failure;
	assert RAM2(2654) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM2(2654))))  severity failure;
	assert RAM2(2655) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM2(2655))))  severity failure;
	assert RAM2(2656) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM2(2656))))  severity failure;
	assert RAM2(2657) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM2(2657))))  severity failure;
	assert RAM2(2658) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM2(2658))))  severity failure;
	assert RAM2(2659) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM2(2659))))  severity failure;
	assert RAM2(2660) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM2(2660))))  severity failure;
	assert RAM2(2661) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM2(2661))))  severity failure;
	assert RAM2(2662) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM2(2662))))  severity failure;
	assert RAM2(2663) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM2(2663))))  severity failure;
	assert RAM2(2664) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM2(2664))))  severity failure;
	assert RAM2(2665) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM2(2665))))  severity failure;
	assert RAM2(2666) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM2(2666))))  severity failure;
	assert RAM2(2667) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM2(2667))))  severity failure;
	assert RAM2(2668) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM2(2668))))  severity failure;
	assert RAM2(2669) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM2(2669))))  severity failure;
	assert RAM2(2670) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM2(2670))))  severity failure;
	assert RAM2(2671) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM2(2671))))  severity failure;
	assert RAM2(2672) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM2(2672))))  severity failure;
	assert RAM2(2673) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM2(2673))))  severity failure;
	assert RAM2(2674) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM2(2674))))  severity failure;
	assert RAM2(2675) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM2(2675))))  severity failure;
	assert RAM2(2676) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM2(2676))))  severity failure;
	assert RAM2(2677) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM2(2677))))  severity failure;
	assert RAM2(2678) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM2(2678))))  severity failure;
	assert RAM2(2679) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM2(2679))))  severity failure;
	assert RAM2(2680) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM2(2680))))  severity failure;
	assert RAM2(2681) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM2(2681))))  severity failure;
	assert RAM2(2682) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM2(2682))))  severity failure;
	assert RAM2(2683) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM2(2683))))  severity failure;
	assert RAM2(2684) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM2(2684))))  severity failure;
	assert RAM2(2685) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM2(2685))))  severity failure;
	assert RAM2(2686) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM2(2686))))  severity failure;
	assert RAM2(2687) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM2(2687))))  severity failure;
	assert RAM2(2688) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM2(2688))))  severity failure;
	assert RAM2(2689) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM2(2689))))  severity failure;
	assert RAM2(2690) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM2(2690))))  severity failure;
	assert RAM2(2691) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM2(2691))))  severity failure;
	assert RAM2(2692) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM2(2692))))  severity failure;
	assert RAM2(2693) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM2(2693))))  severity failure;
	assert RAM2(2694) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM2(2694))))  severity failure;
	assert RAM2(2695) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM2(2695))))  severity failure;
	assert RAM2(2696) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM2(2696))))  severity failure;
	assert RAM2(2697) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM2(2697))))  severity failure;
	assert RAM2(2698) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM2(2698))))  severity failure;
	assert RAM2(2699) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM2(2699))))  severity failure;
	assert RAM2(2700) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM2(2700))))  severity failure;
	assert RAM2(2701) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM2(2701))))  severity failure;
	assert RAM2(2702) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM2(2702))))  severity failure;
	assert RAM2(2703) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM2(2703))))  severity failure;
	assert RAM2(2704) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM2(2704))))  severity failure;
	assert RAM2(2705) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM2(2705))))  severity failure;
	assert RAM2(2706) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM2(2706))))  severity failure;
	assert RAM2(2707) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM2(2707))))  severity failure;
	assert RAM2(2708) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM2(2708))))  severity failure;
	assert RAM2(2709) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM2(2709))))  severity failure;
	assert RAM2(2710) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM2(2710))))  severity failure;
	assert RAM2(2711) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM2(2711))))  severity failure;
	assert RAM2(2712) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM2(2712))))  severity failure;
	assert RAM2(2713) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM2(2713))))  severity failure;
	assert RAM2(2714) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM2(2714))))  severity failure;
	assert RAM2(2715) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM2(2715))))  severity failure;
	assert RAM2(2716) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM2(2716))))  severity failure;
	assert RAM2(2717) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM2(2717))))  severity failure;
	assert RAM2(2718) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM2(2718))))  severity failure;
	assert RAM2(2719) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM2(2719))))  severity failure;
	assert RAM2(2720) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM2(2720))))  severity failure;
	assert RAM2(2721) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM2(2721))))  severity failure;
	assert RAM2(2722) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM2(2722))))  severity failure;
	assert RAM2(2723) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM2(2723))))  severity failure;
	assert RAM2(2724) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM2(2724))))  severity failure;
	assert RAM2(2725) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM2(2725))))  severity failure;
	assert RAM2(2726) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM2(2726))))  severity failure;
	assert RAM2(2727) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM2(2727))))  severity failure;
	assert RAM2(2728) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM2(2728))))  severity failure;
	assert RAM2(2729) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM2(2729))))  severity failure;
	assert RAM2(2730) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM2(2730))))  severity failure;
	assert RAM2(2731) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM2(2731))))  severity failure;
	assert RAM2(2732) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM2(2732))))  severity failure;
	assert RAM2(2733) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM2(2733))))  severity failure;
	assert RAM2(2734) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM2(2734))))  severity failure;
	assert RAM2(2735) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM2(2735))))  severity failure;
	assert RAM2(2736) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM2(2736))))  severity failure;
	assert RAM2(2737) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM2(2737))))  severity failure;
	assert RAM2(2738) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM2(2738))))  severity failure;
	assert RAM2(2739) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM2(2739))))  severity failure;
	assert RAM2(2740) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM2(2740))))  severity failure;
	assert RAM2(2741) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM2(2741))))  severity failure;
	assert RAM2(2742) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM2(2742))))  severity failure;
	assert RAM2(2743) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM2(2743))))  severity failure;
	assert RAM2(2744) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM2(2744))))  severity failure;
	assert RAM2(2745) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM2(2745))))  severity failure;
	assert RAM2(2746) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM2(2746))))  severity failure;
	assert RAM2(2747) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM2(2747))))  severity failure;
	assert RAM2(2748) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM2(2748))))  severity failure;
	assert RAM2(2749) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM2(2749))))  severity failure;
	assert RAM2(2750) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM2(2750))))  severity failure;
	assert RAM2(2751) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM2(2751))))  severity failure;
	assert RAM2(2752) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM2(2752))))  severity failure;
	assert RAM2(2753) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM2(2753))))  severity failure;
	assert RAM2(2754) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM2(2754))))  severity failure;
	assert RAM2(2755) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM2(2755))))  severity failure;
	assert RAM2(2756) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM2(2756))))  severity failure;
	assert RAM2(2757) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM2(2757))))  severity failure;
	assert RAM2(2758) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM2(2758))))  severity failure;
	assert RAM2(2759) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM2(2759))))  severity failure;
	assert RAM2(2760) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM2(2760))))  severity failure;
	assert RAM2(2761) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM2(2761))))  severity failure;
	assert RAM2(2762) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM2(2762))))  severity failure;
	assert RAM2(2763) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM2(2763))))  severity failure;
	assert RAM2(2764) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM2(2764))))  severity failure;
	assert RAM2(2765) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM2(2765))))  severity failure;
	assert RAM2(2766) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM2(2766))))  severity failure;
	assert RAM2(2767) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM2(2767))))  severity failure;
	assert RAM2(2768) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM2(2768))))  severity failure;
	assert RAM2(2769) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM2(2769))))  severity failure;
	assert RAM2(2770) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM2(2770))))  severity failure;
	assert RAM2(2771) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM2(2771))))  severity failure;
	assert RAM2(2772) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM2(2772))))  severity failure;
	assert RAM2(2773) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM2(2773))))  severity failure;
	assert RAM2(2774) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM2(2774))))  severity failure;
	assert RAM2(2775) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM2(2775))))  severity failure;
	assert RAM2(2776) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM2(2776))))  severity failure;
	assert RAM2(2777) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM2(2777))))  severity failure;
	assert RAM2(2778) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM2(2778))))  severity failure;
	assert RAM2(2779) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM2(2779))))  severity failure;
	assert RAM2(2780) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM2(2780))))  severity failure;
	assert RAM2(2781) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM2(2781))))  severity failure;
	assert RAM2(2782) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM2(2782))))  severity failure;
	assert RAM2(2783) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM2(2783))))  severity failure;
	assert RAM2(2784) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM2(2784))))  severity failure;
	assert RAM2(2785) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM2(2785))))  severity failure;
	assert RAM2(2786) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM2(2786))))  severity failure;
	assert RAM2(2787) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM2(2787))))  severity failure;
	assert RAM2(2788) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM2(2788))))  severity failure;
	assert RAM2(2789) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM2(2789))))  severity failure;
	assert RAM2(2790) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM2(2790))))  severity failure;
	assert RAM2(2791) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM2(2791))))  severity failure;
	assert RAM2(2792) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM2(2792))))  severity failure;
	assert RAM2(2793) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM2(2793))))  severity failure;
	assert RAM2(2794) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM2(2794))))  severity failure;
	assert RAM2(2795) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM2(2795))))  severity failure;
	assert RAM2(2796) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM2(2796))))  severity failure;
	assert RAM2(2797) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM2(2797))))  severity failure;
	assert RAM2(2798) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM2(2798))))  severity failure;
	assert RAM2(2799) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM2(2799))))  severity failure;
	assert RAM2(2800) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM2(2800))))  severity failure;
	assert RAM2(2801) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM2(2801))))  severity failure;
	assert RAM2(2802) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM2(2802))))  severity failure;
	assert RAM2(2803) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM2(2803))))  severity failure;
	assert RAM2(2804) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM2(2804))))  severity failure;
	assert RAM2(2805) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM2(2805))))  severity failure;
	assert RAM2(2806) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM2(2806))))  severity failure;
	assert RAM2(2807) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM2(2807))))  severity failure;
	assert RAM2(2808) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM2(2808))))  severity failure;
	assert RAM2(2809) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM2(2809))))  severity failure;
	assert RAM2(2810) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM2(2810))))  severity failure;
	assert RAM2(2811) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM2(2811))))  severity failure;
	assert RAM2(2812) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM2(2812))))  severity failure;
	assert RAM2(2813) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM2(2813))))  severity failure;
	assert RAM2(2814) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM2(2814))))  severity failure;
	assert RAM2(2815) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM2(2815))))  severity failure;
	assert RAM2(2816) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM2(2816))))  severity failure;
	assert RAM2(2817) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM2(2817))))  severity failure;
	assert RAM2(2818) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM2(2818))))  severity failure;
	assert RAM2(2819) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM2(2819))))  severity failure;
	assert RAM2(2820) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM2(2820))))  severity failure;
	assert RAM2(2821) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM2(2821))))  severity failure;
	assert RAM2(2822) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM2(2822))))  severity failure;
	assert RAM2(2823) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM2(2823))))  severity failure;
	assert RAM2(2824) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM2(2824))))  severity failure;
	assert RAM2(2825) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM2(2825))))  severity failure;
	assert RAM2(2826) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM2(2826))))  severity failure;
	assert RAM2(2827) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM2(2827))))  severity failure;
	assert RAM2(2828) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM2(2828))))  severity failure;
	assert RAM2(2829) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM2(2829))))  severity failure;
	assert RAM2(2830) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM2(2830))))  severity failure;
	assert RAM2(2831) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM2(2831))))  severity failure;
	assert RAM2(2832) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM2(2832))))  severity failure;
	assert RAM2(2833) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM2(2833))))  severity failure;
	assert RAM2(2834) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM2(2834))))  severity failure;
	assert RAM2(2835) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM2(2835))))  severity failure;
	assert RAM2(2836) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM2(2836))))  severity failure;
	assert RAM2(2837) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM2(2837))))  severity failure;
	assert RAM2(2838) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM2(2838))))  severity failure;
	assert RAM2(2839) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM2(2839))))  severity failure;
	assert RAM2(2840) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM2(2840))))  severity failure;
	assert RAM2(2841) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM2(2841))))  severity failure;
	assert RAM2(2842) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM2(2842))))  severity failure;
	assert RAM2(2843) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM2(2843))))  severity failure;
	assert RAM2(2844) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM2(2844))))  severity failure;
	assert RAM2(2845) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM2(2845))))  severity failure;
	assert RAM2(2846) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM2(2846))))  severity failure;
	assert RAM2(2847) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM2(2847))))  severity failure;
	assert RAM2(2848) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM2(2848))))  severity failure;
	assert RAM2(2849) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM2(2849))))  severity failure;
	assert RAM2(2850) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM2(2850))))  severity failure;
	assert RAM2(2851) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM2(2851))))  severity failure;
	assert RAM2(2852) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM2(2852))))  severity failure;
	assert RAM2(2853) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM2(2853))))  severity failure;
	assert RAM2(2854) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM2(2854))))  severity failure;
	assert RAM2(2855) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM2(2855))))  severity failure;
	assert RAM2(2856) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM2(2856))))  severity failure;
	assert RAM2(2857) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM2(2857))))  severity failure;
	assert RAM2(2858) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM2(2858))))  severity failure;
	assert RAM2(2859) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM2(2859))))  severity failure;
	assert RAM2(2860) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM2(2860))))  severity failure;
	assert RAM2(2861) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM2(2861))))  severity failure;
	assert RAM2(2862) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM2(2862))))  severity failure;
	assert RAM2(2863) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM2(2863))))  severity failure;
	assert RAM2(2864) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM2(2864))))  severity failure;
	assert RAM2(2865) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM2(2865))))  severity failure;
	assert RAM2(2866) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM2(2866))))  severity failure;
	assert RAM2(2867) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM2(2867))))  severity failure;
	assert RAM2(2868) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM2(2868))))  severity failure;
	assert RAM2(2869) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM2(2869))))  severity failure;
	assert RAM2(2870) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM2(2870))))  severity failure;
	assert RAM2(2871) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM2(2871))))  severity failure;
	assert RAM2(2872) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM2(2872))))  severity failure;
	assert RAM2(2873) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM2(2873))))  severity failure;
	assert RAM2(2874) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM2(2874))))  severity failure;
	assert RAM2(2875) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM2(2875))))  severity failure;
	assert RAM2(2876) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM2(2876))))  severity failure;
	assert RAM2(2877) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM2(2877))))  severity failure;
	assert RAM2(2878) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM2(2878))))  severity failure;
	assert RAM2(2879) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM2(2879))))  severity failure;
	assert RAM2(2880) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM2(2880))))  severity failure;
	assert RAM2(2881) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM2(2881))))  severity failure;
	assert RAM2(2882) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM2(2882))))  severity failure;
	assert RAM2(2883) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM2(2883))))  severity failure;
	assert RAM2(2884) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM2(2884))))  severity failure;
	assert RAM2(2885) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM2(2885))))  severity failure;
	assert RAM2(2886) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM2(2886))))  severity failure;
	assert RAM2(2887) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM2(2887))))  severity failure;
	assert RAM2(2888) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM2(2888))))  severity failure;
	assert RAM2(2889) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM2(2889))))  severity failure;
	assert RAM2(2890) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM2(2890))))  severity failure;
	assert RAM2(2891) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM2(2891))))  severity failure;
	assert RAM2(2892) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM2(2892))))  severity failure;
	assert RAM2(2893) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM2(2893))))  severity failure;
	assert RAM2(2894) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM2(2894))))  severity failure;
	assert RAM2(2895) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM2(2895))))  severity failure;
	assert RAM2(2896) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM2(2896))))  severity failure;
	assert RAM2(2897) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM2(2897))))  severity failure;
	assert RAM2(2898) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM2(2898))))  severity failure;
	assert RAM2(2899) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM2(2899))))  severity failure;
	assert RAM2(2900) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM2(2900))))  severity failure;
	assert RAM2(2901) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM2(2901))))  severity failure;
	assert RAM2(2902) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM2(2902))))  severity failure;
	assert RAM2(2903) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM2(2903))))  severity failure;
	assert RAM2(2904) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM2(2904))))  severity failure;
	assert RAM2(2905) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM2(2905))))  severity failure;
	assert RAM2(2906) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM2(2906))))  severity failure;
	assert RAM2(2907) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM2(2907))))  severity failure;
	assert RAM2(2908) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM2(2908))))  severity failure;
	assert RAM2(2909) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM2(2909))))  severity failure;
	assert RAM2(2910) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM2(2910))))  severity failure;
	assert RAM2(2911) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM2(2911))))  severity failure;
	assert RAM2(2912) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM2(2912))))  severity failure;
	assert RAM2(2913) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM2(2913))))  severity failure;
	assert RAM2(2914) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM2(2914))))  severity failure;
	assert RAM2(2915) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM2(2915))))  severity failure;
	assert RAM2(2916) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM2(2916))))  severity failure;
	assert RAM2(2917) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM2(2917))))  severity failure;
	assert RAM2(2918) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM2(2918))))  severity failure;
	assert RAM2(2919) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM2(2919))))  severity failure;
	assert RAM2(2920) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM2(2920))))  severity failure;
	assert RAM2(2921) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM2(2921))))  severity failure;
	assert RAM2(2922) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM2(2922))))  severity failure;
	assert RAM2(2923) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM2(2923))))  severity failure;
	assert RAM2(2924) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM2(2924))))  severity failure;
	assert RAM2(2925) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM2(2925))))  severity failure;
	assert RAM2(2926) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM2(2926))))  severity failure;
	assert RAM2(2927) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM2(2927))))  severity failure;
	assert RAM2(2928) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM2(2928))))  severity failure;
	assert RAM2(2929) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM2(2929))))  severity failure;
	assert RAM2(2930) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM2(2930))))  severity failure;
	assert RAM2(2931) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM2(2931))))  severity failure;
	assert RAM2(2932) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM2(2932))))  severity failure;
	assert RAM2(2933) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM2(2933))))  severity failure;
	assert RAM2(2934) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM2(2934))))  severity failure;
	assert RAM2(2935) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM2(2935))))  severity failure;
	assert RAM2(2936) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM2(2936))))  severity failure;
	assert RAM2(2937) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM2(2937))))  severity failure;
	assert RAM2(2938) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM2(2938))))  severity failure;
	assert RAM2(2939) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM2(2939))))  severity failure;
	assert RAM2(2940) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM2(2940))))  severity failure;
	assert RAM2(2941) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM2(2941))))  severity failure;
	assert RAM2(2942) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM2(2942))))  severity failure;
	assert RAM2(2943) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM2(2943))))  severity failure;
	assert RAM2(2944) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM2(2944))))  severity failure;
	assert RAM2(2945) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM2(2945))))  severity failure;
	assert RAM2(2946) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM2(2946))))  severity failure;
	assert RAM2(2947) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM2(2947))))  severity failure;
	assert RAM2(2948) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM2(2948))))  severity failure;
	assert RAM2(2949) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM2(2949))))  severity failure;
	assert RAM2(2950) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM2(2950))))  severity failure;
	assert RAM2(2951) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM2(2951))))  severity failure;
	assert RAM2(2952) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM2(2952))))  severity failure;
	assert RAM2(2953) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM2(2953))))  severity failure;
	assert RAM2(2954) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM2(2954))))  severity failure;
	assert RAM2(2955) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM2(2955))))  severity failure;
	assert RAM2(2956) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM2(2956))))  severity failure;
	assert RAM2(2957) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM2(2957))))  severity failure;
	assert RAM2(2958) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM2(2958))))  severity failure;
	assert RAM2(2959) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM2(2959))))  severity failure;
	assert RAM2(2960) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM2(2960))))  severity failure;
	assert RAM2(2961) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM2(2961))))  severity failure;
	assert RAM2(2962) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM2(2962))))  severity failure;
	assert RAM2(2963) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM2(2963))))  severity failure;
	assert RAM2(2964) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM2(2964))))  severity failure;
	assert RAM2(2965) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM2(2965))))  severity failure;
	assert RAM2(2966) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM2(2966))))  severity failure;
	assert RAM2(2967) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM2(2967))))  severity failure;
	assert RAM2(2968) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM2(2968))))  severity failure;
	assert RAM2(2969) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM2(2969))))  severity failure;
	assert RAM2(2970) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM2(2970))))  severity failure;
	assert RAM2(2971) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM2(2971))))  severity failure;
	assert RAM2(2972) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM2(2972))))  severity failure;
	assert RAM2(2973) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM2(2973))))  severity failure;
	assert RAM2(2974) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM2(2974))))  severity failure;
	assert RAM2(2975) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM2(2975))))  severity failure;
	assert RAM2(2976) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM2(2976))))  severity failure;
	assert RAM2(2977) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM2(2977))))  severity failure;
	assert RAM2(2978) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM2(2978))))  severity failure;
	assert RAM2(2979) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM2(2979))))  severity failure;
	assert RAM2(2980) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM2(2980))))  severity failure;
	assert RAM2(2981) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM2(2981))))  severity failure;
	assert RAM2(2982) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM2(2982))))  severity failure;
	assert RAM2(2983) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM2(2983))))  severity failure;
	assert RAM2(2984) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM2(2984))))  severity failure;
	assert RAM2(2985) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM2(2985))))  severity failure;
	assert RAM2(2986) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM2(2986))))  severity failure;
	assert RAM2(2987) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM2(2987))))  severity failure;
	assert RAM2(2988) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM2(2988))))  severity failure;
	assert RAM2(2989) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM2(2989))))  severity failure;
	assert RAM2(2990) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM2(2990))))  severity failure;
	assert RAM2(2991) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM2(2991))))  severity failure;
	assert RAM2(2992) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM2(2992))))  severity failure;
	assert RAM2(2993) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM2(2993))))  severity failure;
	assert RAM2(2994) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM2(2994))))  severity failure;
	assert RAM2(2995) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM2(2995))))  severity failure;
	assert RAM2(2996) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM2(2996))))  severity failure;
	assert RAM2(2997) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM2(2997))))  severity failure;
	assert RAM2(2998) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM2(2998))))  severity failure;
	assert RAM2(2999) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM2(2999))))  severity failure;
	assert RAM2(3000) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM2(3000))))  severity failure;
	assert RAM2(3001) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM2(3001))))  severity failure;
	assert RAM2(3002) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM2(3002))))  severity failure;
	assert RAM2(3003) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM2(3003))))  severity failure;
	assert RAM2(3004) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM2(3004))))  severity failure;
	assert RAM2(3005) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM2(3005))))  severity failure;
	assert RAM2(3006) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM2(3006))))  severity failure;
	assert RAM2(3007) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM2(3007))))  severity failure;
	assert RAM2(3008) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM2(3008))))  severity failure;
	assert RAM2(3009) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM2(3009))))  severity failure;
	assert RAM2(3010) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM2(3010))))  severity failure;
	assert RAM2(3011) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM2(3011))))  severity failure;
	assert RAM2(3012) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM2(3012))))  severity failure;
	assert RAM2(3013) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM2(3013))))  severity failure;
	assert RAM2(3014) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM2(3014))))  severity failure;
	assert RAM2(3015) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM2(3015))))  severity failure;
	assert RAM2(3016) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM2(3016))))  severity failure;
	assert RAM2(3017) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM2(3017))))  severity failure;
	assert RAM2(3018) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM2(3018))))  severity failure;
	assert RAM2(3019) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM2(3019))))  severity failure;
	assert RAM2(3020) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM2(3020))))  severity failure;
	assert RAM2(3021) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM2(3021))))  severity failure;
	assert RAM2(3022) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM2(3022))))  severity failure;
	assert RAM2(3023) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM2(3023))))  severity failure;
	assert RAM2(3024) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM2(3024))))  severity failure;
	assert RAM2(3025) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM2(3025))))  severity failure;
	assert RAM2(3026) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM2(3026))))  severity failure;
	assert RAM2(3027) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM2(3027))))  severity failure;
	assert RAM2(3028) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM2(3028))))  severity failure;
	assert RAM2(3029) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM2(3029))))  severity failure;
	assert RAM2(3030) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM2(3030))))  severity failure;
	assert RAM2(3031) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM2(3031))))  severity failure;
	assert RAM2(3032) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM2(3032))))  severity failure;
	assert RAM2(3033) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM2(3033))))  severity failure;
	assert RAM2(3034) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM2(3034))))  severity failure;
	assert RAM2(3035) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM2(3035))))  severity failure;
	assert RAM2(3036) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM2(3036))))  severity failure;
	assert RAM2(3037) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM2(3037))))  severity failure;
	assert RAM2(3038) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM2(3038))))  severity failure;
	assert RAM2(3039) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM2(3039))))  severity failure;
	assert RAM2(3040) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM2(3040))))  severity failure;
	assert RAM2(3041) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM2(3041))))  severity failure;
	assert RAM2(3042) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM2(3042))))  severity failure;
	assert RAM2(3043) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM2(3043))))  severity failure;
	assert RAM2(3044) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM2(3044))))  severity failure;
	assert RAM2(3045) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM2(3045))))  severity failure;
	assert RAM2(3046) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM2(3046))))  severity failure;
	assert RAM2(3047) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM2(3047))))  severity failure;
	assert RAM2(3048) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM2(3048))))  severity failure;
	assert RAM2(3049) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM2(3049))))  severity failure;
	assert RAM2(3050) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM2(3050))))  severity failure;
	assert RAM2(3051) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM2(3051))))  severity failure;
	assert RAM2(3052) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM2(3052))))  severity failure;
	assert RAM2(3053) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM2(3053))))  severity failure;
	assert RAM2(3054) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM2(3054))))  severity failure;
	assert RAM2(3055) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM2(3055))))  severity failure;
	assert RAM2(3056) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM2(3056))))  severity failure;
	assert RAM2(3057) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM2(3057))))  severity failure;
	assert RAM2(3058) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM2(3058))))  severity failure;
	assert RAM2(3059) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM2(3059))))  severity failure;
	assert RAM2(3060) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM2(3060))))  severity failure;
	assert RAM2(3061) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM2(3061))))  severity failure;
	assert RAM2(3062) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM2(3062))))  severity failure;
	assert RAM2(3063) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM2(3063))))  severity failure;
	assert RAM2(3064) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM2(3064))))  severity failure;
	assert RAM2(3065) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM2(3065))))  severity failure;
	assert RAM2(3066) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM2(3066))))  severity failure;
	assert RAM2(3067) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM2(3067))))  severity failure;
	assert RAM2(3068) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM2(3068))))  severity failure;
	assert RAM2(3069) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM2(3069))))  severity failure;
	assert RAM2(3070) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM2(3070))))  severity failure;
	assert RAM2(3071) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM2(3071))))  severity failure;
	assert RAM2(3072) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM2(3072))))  severity failure;
	assert RAM2(3073) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM2(3073))))  severity failure;
	assert RAM2(3074) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM2(3074))))  severity failure;
	assert RAM2(3075) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM2(3075))))  severity failure;
	assert RAM2(3076) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM2(3076))))  severity failure;
	assert RAM2(3077) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM2(3077))))  severity failure;
	assert RAM2(3078) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM2(3078))))  severity failure;
	assert RAM2(3079) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM2(3079))))  severity failure;
	assert RAM2(3080) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM2(3080))))  severity failure;
	assert RAM2(3081) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM2(3081))))  severity failure;
	assert RAM2(3082) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM2(3082))))  severity failure;
	assert RAM2(3083) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM2(3083))))  severity failure;
	assert RAM2(3084) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM2(3084))))  severity failure;
	assert RAM2(3085) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM2(3085))))  severity failure;
	assert RAM2(3086) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM2(3086))))  severity failure;
	assert RAM2(3087) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM2(3087))))  severity failure;
	assert RAM2(3088) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM2(3088))))  severity failure;
	assert RAM2(3089) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM2(3089))))  severity failure;
	assert RAM2(3090) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM2(3090))))  severity failure;
	assert RAM2(3091) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM2(3091))))  severity failure;
	assert RAM2(3092) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM2(3092))))  severity failure;
	assert RAM2(3093) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM2(3093))))  severity failure;
	assert RAM2(3094) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM2(3094))))  severity failure;
	assert RAM2(3095) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM2(3095))))  severity failure;
	assert RAM2(3096) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM2(3096))))  severity failure;
	assert RAM2(3097) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM2(3097))))  severity failure;
	assert RAM2(3098) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM2(3098))))  severity failure;
	assert RAM2(3099) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM2(3099))))  severity failure;
	assert RAM2(3100) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM2(3100))))  severity failure;
	assert RAM2(3101) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM2(3101))))  severity failure;
	assert RAM2(3102) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM2(3102))))  severity failure;
	assert RAM2(3103) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM2(3103))))  severity failure;
	assert RAM2(3104) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM2(3104))))  severity failure;
	assert RAM2(3105) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM2(3105))))  severity failure;
	assert RAM2(3106) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM2(3106))))  severity failure;
	assert RAM2(3107) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM2(3107))))  severity failure;
	assert RAM2(3108) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM2(3108))))  severity failure;
	assert RAM2(3109) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM2(3109))))  severity failure;
	assert RAM2(3110) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM2(3110))))  severity failure;
	assert RAM2(3111) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM2(3111))))  severity failure;
	assert RAM2(3112) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM2(3112))))  severity failure;
	assert RAM2(3113) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM2(3113))))  severity failure;
	assert RAM2(3114) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM2(3114))))  severity failure;
	assert RAM2(3115) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM2(3115))))  severity failure;
	assert RAM2(3116) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM2(3116))))  severity failure;
	assert RAM2(3117) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM2(3117))))  severity failure;
	assert RAM2(3118) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM2(3118))))  severity failure;
	assert RAM2(3119) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM2(3119))))  severity failure;
	assert RAM2(3120) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM2(3120))))  severity failure;
	assert RAM2(3121) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM2(3121))))  severity failure;
	assert RAM2(3122) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM2(3122))))  severity failure;
	assert RAM2(3123) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM2(3123))))  severity failure;
	assert RAM2(3124) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM2(3124))))  severity failure;
	assert RAM2(3125) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM2(3125))))  severity failure;
	assert RAM2(3126) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM2(3126))))  severity failure;
	assert RAM2(3127) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM2(3127))))  severity failure;
	assert RAM2(3128) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM2(3128))))  severity failure;
	assert RAM2(3129) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM2(3129))))  severity failure;
	assert RAM2(3130) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM2(3130))))  severity failure;
	assert RAM2(3131) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM2(3131))))  severity failure;
	assert RAM2(3132) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM2(3132))))  severity failure;
	assert RAM2(3133) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM2(3133))))  severity failure;
	assert RAM2(3134) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM2(3134))))  severity failure;
	assert RAM2(3135) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM2(3135))))  severity failure;
	assert RAM2(3136) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM2(3136))))  severity failure;
	assert RAM2(3137) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM2(3137))))  severity failure;
	assert RAM2(3138) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM2(3138))))  severity failure;
	assert RAM2(3139) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM2(3139))))  severity failure;
	assert RAM2(3140) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM2(3140))))  severity failure;
	assert RAM2(3141) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM2(3141))))  severity failure;
	assert RAM2(3142) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM2(3142))))  severity failure;
	assert RAM2(3143) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM2(3143))))  severity failure;
	assert RAM2(3144) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM2(3144))))  severity failure;
	assert RAM2(3145) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM2(3145))))  severity failure;
	assert RAM2(3146) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM2(3146))))  severity failure;
	assert RAM2(3147) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM2(3147))))  severity failure;
	assert RAM2(3148) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM2(3148))))  severity failure;
	assert RAM2(3149) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM2(3149))))  severity failure;
	assert RAM2(3150) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM2(3150))))  severity failure;
	assert RAM2(3151) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM2(3151))))  severity failure;
	assert RAM2(3152) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM2(3152))))  severity failure;
	assert RAM2(3153) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM2(3153))))  severity failure;
	assert RAM2(3154) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM2(3154))))  severity failure;
	assert RAM2(3155) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM2(3155))))  severity failure;
	assert RAM2(3156) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM2(3156))))  severity failure;
	assert RAM2(3157) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM2(3157))))  severity failure;
	assert RAM2(3158) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM2(3158))))  severity failure;
	assert RAM2(3159) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM2(3159))))  severity failure;
	assert RAM2(3160) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM2(3160))))  severity failure;
	assert RAM2(3161) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM2(3161))))  severity failure;
	assert RAM2(3162) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM2(3162))))  severity failure;
	assert RAM2(3163) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM2(3163))))  severity failure;
	assert RAM2(3164) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM2(3164))))  severity failure;
	assert RAM2(3165) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM2(3165))))  severity failure;
	assert RAM2(3166) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM2(3166))))  severity failure;
	assert RAM2(3167) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM2(3167))))  severity failure;
	assert RAM2(3168) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM2(3168))))  severity failure;
	assert RAM2(3169) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM2(3169))))  severity failure;
	assert RAM2(3170) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM2(3170))))  severity failure;
	assert RAM2(3171) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM2(3171))))  severity failure;
	assert RAM2(3172) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM2(3172))))  severity failure;
	assert RAM2(3173) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM2(3173))))  severity failure;
	assert RAM2(3174) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM2(3174))))  severity failure;
	assert RAM2(3175) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM2(3175))))  severity failure;
	assert RAM2(3176) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM2(3176))))  severity failure;
	assert RAM2(3177) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM2(3177))))  severity failure;
	assert RAM2(3178) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM2(3178))))  severity failure;
	assert RAM2(3179) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM2(3179))))  severity failure;
	assert RAM2(3180) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM2(3180))))  severity failure;
	assert RAM2(3181) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM2(3181))))  severity failure;
	assert RAM2(3182) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM2(3182))))  severity failure;
	assert RAM2(3183) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM2(3183))))  severity failure;
	assert RAM2(3184) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM2(3184))))  severity failure;
	assert RAM2(3185) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM2(3185))))  severity failure;
	assert RAM2(3186) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM2(3186))))  severity failure;
	assert RAM2(3187) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM2(3187))))  severity failure;
	assert RAM2(3188) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM2(3188))))  severity failure;
	assert RAM2(3189) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM2(3189))))  severity failure;
	assert RAM2(3190) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM2(3190))))  severity failure;
	assert RAM2(3191) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM2(3191))))  severity failure;
	assert RAM2(3192) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM2(3192))))  severity failure;
	assert RAM2(3193) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM2(3193))))  severity failure;
	assert RAM2(3194) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM2(3194))))  severity failure;
	assert RAM2(3195) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM2(3195))))  severity failure;
	assert RAM2(3196) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM2(3196))))  severity failure;
	assert RAM2(3197) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM2(3197))))  severity failure;
	assert RAM2(3198) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM2(3198))))  severity failure;
	assert RAM2(3199) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM2(3199))))  severity failure;
	assert RAM2(3200) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM2(3200))))  severity failure;
	assert RAM2(3201) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM2(3201))))  severity failure;
	assert RAM2(3202) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM2(3202))))  severity failure;
	assert RAM2(3203) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM2(3203))))  severity failure;
	assert RAM2(3204) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM2(3204))))  severity failure;
	assert RAM2(3205) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM2(3205))))  severity failure;
	assert RAM2(3206) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM2(3206))))  severity failure;
	assert RAM2(3207) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM2(3207))))  severity failure;
	assert RAM2(3208) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM2(3208))))  severity failure;
	assert RAM2(3209) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM2(3209))))  severity failure;
	assert RAM2(3210) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM2(3210))))  severity failure;
	assert RAM2(3211) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM2(3211))))  severity failure;
	assert RAM2(3212) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM2(3212))))  severity failure;
	assert RAM2(3213) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM2(3213))))  severity failure;
	assert RAM2(3214) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM2(3214))))  severity failure;
	assert RAM2(3215) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM2(3215))))  severity failure;
	assert RAM2(3216) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM2(3216))))  severity failure;
	assert RAM2(3217) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM2(3217))))  severity failure;
	assert RAM2(3218) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM2(3218))))  severity failure;
	assert RAM2(3219) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM2(3219))))  severity failure;
	assert RAM2(3220) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM2(3220))))  severity failure;
	assert RAM2(3221) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM2(3221))))  severity failure;
	assert RAM2(3222) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM2(3222))))  severity failure;
	assert RAM2(3223) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM2(3223))))  severity failure;
	assert RAM2(3224) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM2(3224))))  severity failure;
	assert RAM2(3225) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM2(3225))))  severity failure;
	assert RAM2(3226) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM2(3226))))  severity failure;
	assert RAM2(3227) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM2(3227))))  severity failure;
	assert RAM2(3228) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM2(3228))))  severity failure;
	assert RAM2(3229) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM2(3229))))  severity failure;
	assert RAM2(3230) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM2(3230))))  severity failure;
	assert RAM2(3231) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM2(3231))))  severity failure;
	assert RAM2(3232) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM2(3232))))  severity failure;
	assert RAM2(3233) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM2(3233))))  severity failure;
	assert RAM2(3234) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM2(3234))))  severity failure;
	assert RAM2(3235) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM2(3235))))  severity failure;
	assert RAM2(3236) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM2(3236))))  severity failure;
	assert RAM2(3237) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM2(3237))))  severity failure;
	assert RAM2(3238) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM2(3238))))  severity failure;
	assert RAM2(3239) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM2(3239))))  severity failure;
	assert RAM2(3240) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM2(3240))))  severity failure;
	assert RAM2(3241) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM2(3241))))  severity failure;
	assert RAM2(3242) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM2(3242))))  severity failure;
	assert RAM2(3243) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM2(3243))))  severity failure;
	assert RAM2(3244) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM2(3244))))  severity failure;
	assert RAM2(3245) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM2(3245))))  severity failure;
	assert RAM2(3246) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM2(3246))))  severity failure;
	assert RAM2(3247) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM2(3247))))  severity failure;
	assert RAM2(3248) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM2(3248))))  severity failure;
	assert RAM2(3249) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM2(3249))))  severity failure;
	assert RAM2(3250) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM2(3250))))  severity failure;
	assert RAM2(3251) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM2(3251))))  severity failure;
	assert RAM2(3252) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM2(3252))))  severity failure;
	assert RAM2(3253) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM2(3253))))  severity failure;
	assert RAM2(3254) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM2(3254))))  severity failure;
	assert RAM2(3255) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM2(3255))))  severity failure;
	assert RAM2(3256) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM2(3256))))  severity failure;
	assert RAM2(3257) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM2(3257))))  severity failure;
	assert RAM2(3258) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM2(3258))))  severity failure;
	assert RAM2(3259) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM2(3259))))  severity failure;
	assert RAM2(3260) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM2(3260))))  severity failure;
	assert RAM2(3261) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM2(3261))))  severity failure;
	assert RAM2(3262) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM2(3262))))  severity failure;
	assert RAM2(3263) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM2(3263))))  severity failure;
	assert RAM2(3264) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM2(3264))))  severity failure;
	assert RAM2(3265) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM2(3265))))  severity failure;
	assert RAM2(3266) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM2(3266))))  severity failure;
	assert RAM2(3267) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM2(3267))))  severity failure;
	assert RAM2(3268) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM2(3268))))  severity failure;
	assert RAM2(3269) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM2(3269))))  severity failure;
	assert RAM2(3270) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM2(3270))))  severity failure;
	assert RAM2(3271) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM2(3271))))  severity failure;
	assert RAM2(3272) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM2(3272))))  severity failure;
	assert RAM2(3273) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM2(3273))))  severity failure;
	assert RAM2(3274) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM2(3274))))  severity failure;
	assert RAM2(3275) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM2(3275))))  severity failure;
	assert RAM2(3276) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM2(3276))))  severity failure;
	assert RAM2(3277) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM2(3277))))  severity failure;
	assert RAM2(3278) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM2(3278))))  severity failure;
	assert RAM2(3279) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM2(3279))))  severity failure;
	assert RAM2(3280) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM2(3280))))  severity failure;
	assert RAM2(3281) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM2(3281))))  severity failure;
	assert RAM2(3282) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM2(3282))))  severity failure;
	assert RAM2(3283) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM2(3283))))  severity failure;
	assert RAM2(3284) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM2(3284))))  severity failure;
	assert RAM2(3285) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM2(3285))))  severity failure;
	assert RAM2(3286) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM2(3286))))  severity failure;
	assert RAM2(3287) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM2(3287))))  severity failure;
	assert RAM2(3288) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM2(3288))))  severity failure;
	assert RAM2(3289) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM2(3289))))  severity failure;
	assert RAM2(3290) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM2(3290))))  severity failure;
	assert RAM2(3291) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM2(3291))))  severity failure;
	assert RAM2(3292) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM2(3292))))  severity failure;
	assert RAM2(3293) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM2(3293))))  severity failure;
	assert RAM2(3294) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM2(3294))))  severity failure;
	assert RAM2(3295) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM2(3295))))  severity failure;
	assert RAM2(3296) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM2(3296))))  severity failure;
	assert RAM2(3297) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM2(3297))))  severity failure;
	assert RAM2(3298) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM2(3298))))  severity failure;
	assert RAM2(3299) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM2(3299))))  severity failure;
	assert RAM2(3300) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM2(3300))))  severity failure;
	assert RAM2(3301) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM2(3301))))  severity failure;
	assert RAM2(3302) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM2(3302))))  severity failure;
	assert RAM2(3303) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM2(3303))))  severity failure;
	assert RAM2(3304) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM2(3304))))  severity failure;
	assert RAM2(3305) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM2(3305))))  severity failure;
	assert RAM2(3306) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM2(3306))))  severity failure;
	assert RAM2(3307) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM2(3307))))  severity failure;
	assert RAM2(3308) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM2(3308))))  severity failure;
	assert RAM2(3309) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM2(3309))))  severity failure;
	assert RAM2(3310) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM2(3310))))  severity failure;
	assert RAM2(3311) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM2(3311))))  severity failure;
	assert RAM2(3312) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM2(3312))))  severity failure;
	assert RAM2(3313) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM2(3313))))  severity failure;


    assert false report "Simulation Ended! TEST PASSATO" severity failure;
end process test;

end projecttb; 


