
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity project_tb is
end project_tb;

architecture projecttb of project_tb is
constant c_CLOCK_PERIOD         : time := 15 ns;
signal   tb_done                : std_logic;
signal   mem_address            : std_logic_vector (15 downto 0) := (others => '0');
signal   tb_rst                 : std_logic := '0';
signal   tb_start               : std_logic := '0';
signal   tb_clk                 : std_logic := '0';
signal   mem_o_data,mem_i_data  : std_logic_vector (7 downto 0);
signal   enable_wire            : std_logic;
signal   mem_we                 : std_logic;

type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);


signal RAM: ram_type := (
			0 => std_logic_vector(to_unsigned(58, 8)),
			1 => std_logic_vector(to_unsigned(11, 8)),
			2 => std_logic_vector(to_unsigned(164, 8)),
			3 => std_logic_vector(to_unsigned(118, 8)),
			4 => std_logic_vector(to_unsigned(240, 8)),
			5 => std_logic_vector(to_unsigned(22, 8)),
			6 => std_logic_vector(to_unsigned(78, 8)),
			7 => std_logic_vector(to_unsigned(115, 8)),
			8 => std_logic_vector(to_unsigned(41, 8)),
			9 => std_logic_vector(to_unsigned(116, 8)),
			10 => std_logic_vector(to_unsigned(241, 8)),
			11 => std_logic_vector(to_unsigned(43, 8)),
			12 => std_logic_vector(to_unsigned(30, 8)),
			13 => std_logic_vector(to_unsigned(244, 8)),
			14 => std_logic_vector(to_unsigned(45, 8)),
			15 => std_logic_vector(to_unsigned(252, 8)),
			16 => std_logic_vector(to_unsigned(50, 8)),
			17 => std_logic_vector(to_unsigned(134, 8)),
			18 => std_logic_vector(to_unsigned(23, 8)),
			19 => std_logic_vector(to_unsigned(61, 8)),
			20 => std_logic_vector(to_unsigned(205, 8)),
			21 => std_logic_vector(to_unsigned(250, 8)),
			22 => std_logic_vector(to_unsigned(47, 8)),
			23 => std_logic_vector(to_unsigned(120, 8)),
			24 => std_logic_vector(to_unsigned(104, 8)),
			25 => std_logic_vector(to_unsigned(18, 8)),
			26 => std_logic_vector(to_unsigned(53, 8)),
			27 => std_logic_vector(to_unsigned(203, 8)),
			28 => std_logic_vector(to_unsigned(34, 8)),
			29 => std_logic_vector(to_unsigned(192, 8)),
			30 => std_logic_vector(to_unsigned(53, 8)),
			31 => std_logic_vector(to_unsigned(50, 8)),
			32 => std_logic_vector(to_unsigned(27, 8)),
			33 => std_logic_vector(to_unsigned(220, 8)),
			34 => std_logic_vector(to_unsigned(158, 8)),
			35 => std_logic_vector(to_unsigned(7, 8)),
			36 => std_logic_vector(to_unsigned(132, 8)),
			37 => std_logic_vector(to_unsigned(90, 8)),
			38 => std_logic_vector(to_unsigned(216, 8)),
			39 => std_logic_vector(to_unsigned(8, 8)),
			40 => std_logic_vector(to_unsigned(198, 8)),
			41 => std_logic_vector(to_unsigned(159, 8)),
			42 => std_logic_vector(to_unsigned(116, 8)),
			43 => std_logic_vector(to_unsigned(23, 8)),
			44 => std_logic_vector(to_unsigned(157, 8)),
			45 => std_logic_vector(to_unsigned(240, 8)),
			46 => std_logic_vector(to_unsigned(162, 8)),
			47 => std_logic_vector(to_unsigned(225, 8)),
			48 => std_logic_vector(to_unsigned(228, 8)),
			49 => std_logic_vector(to_unsigned(176, 8)),
			50 => std_logic_vector(to_unsigned(161, 8)),
			51 => std_logic_vector(to_unsigned(247, 8)),
			52 => std_logic_vector(to_unsigned(174, 8)),
			53 => std_logic_vector(to_unsigned(223, 8)),
			54 => std_logic_vector(to_unsigned(72, 8)),
			55 => std_logic_vector(to_unsigned(104, 8)),
			56 => std_logic_vector(to_unsigned(91, 8)),
			57 => std_logic_vector(to_unsigned(79, 8)),
			58 => std_logic_vector(to_unsigned(154, 8)),
			59 => std_logic_vector(to_unsigned(126, 8)),
			60 => std_logic_vector(to_unsigned(45, 8)),
			61 => std_logic_vector(to_unsigned(2, 8)),
			62 => std_logic_vector(to_unsigned(116, 8)),
			63 => std_logic_vector(to_unsigned(85, 8)),
			64 => std_logic_vector(to_unsigned(245, 8)),
			65 => std_logic_vector(to_unsigned(26, 8)),
			66 => std_logic_vector(to_unsigned(236, 8)),
			67 => std_logic_vector(to_unsigned(153, 8)),
			68 => std_logic_vector(to_unsigned(100, 8)),
			69 => std_logic_vector(to_unsigned(110, 8)),
			70 => std_logic_vector(to_unsigned(163, 8)),
			71 => std_logic_vector(to_unsigned(227, 8)),
			72 => std_logic_vector(to_unsigned(111, 8)),
			73 => std_logic_vector(to_unsigned(152, 8)),
			74 => std_logic_vector(to_unsigned(0, 8)),
			75 => std_logic_vector(to_unsigned(151, 8)),
			76 => std_logic_vector(to_unsigned(55, 8)),
			77 => std_logic_vector(to_unsigned(36, 8)),
			78 => std_logic_vector(to_unsigned(199, 8)),
			79 => std_logic_vector(to_unsigned(123, 8)),
			80 => std_logic_vector(to_unsigned(73, 8)),
			81 => std_logic_vector(to_unsigned(32, 8)),
			82 => std_logic_vector(to_unsigned(106, 8)),
			83 => std_logic_vector(to_unsigned(40, 8)),
			84 => std_logic_vector(to_unsigned(1, 8)),
			85 => std_logic_vector(to_unsigned(35, 8)),
			86 => std_logic_vector(to_unsigned(121, 8)),
			87 => std_logic_vector(to_unsigned(152, 8)),
			88 => std_logic_vector(to_unsigned(87, 8)),
			89 => std_logic_vector(to_unsigned(27, 8)),
			90 => std_logic_vector(to_unsigned(29, 8)),
			91 => std_logic_vector(to_unsigned(137, 8)),
			92 => std_logic_vector(to_unsigned(232, 8)),
			93 => std_logic_vector(to_unsigned(122, 8)),
			94 => std_logic_vector(to_unsigned(59, 8)),
			95 => std_logic_vector(to_unsigned(12, 8)),
			96 => std_logic_vector(to_unsigned(8, 8)),
			97 => std_logic_vector(to_unsigned(25, 8)),
			98 => std_logic_vector(to_unsigned(6, 8)),
			99 => std_logic_vector(to_unsigned(254, 8)),
			100 => std_logic_vector(to_unsigned(223, 8)),
			101 => std_logic_vector(to_unsigned(21, 8)),
			102 => std_logic_vector(to_unsigned(21, 8)),
			103 => std_logic_vector(to_unsigned(132, 8)),
			104 => std_logic_vector(to_unsigned(174, 8)),
			105 => std_logic_vector(to_unsigned(248, 8)),
			106 => std_logic_vector(to_unsigned(135, 8)),
			107 => std_logic_vector(to_unsigned(236, 8)),
			108 => std_logic_vector(to_unsigned(164, 8)),
			109 => std_logic_vector(to_unsigned(139, 8)),
			110 => std_logic_vector(to_unsigned(64, 8)),
			111 => std_logic_vector(to_unsigned(196, 8)),
			112 => std_logic_vector(to_unsigned(90, 8)),
			113 => std_logic_vector(to_unsigned(45, 8)),
			114 => std_logic_vector(to_unsigned(133, 8)),
			115 => std_logic_vector(to_unsigned(210, 8)),
			116 => std_logic_vector(to_unsigned(115, 8)),
			117 => std_logic_vector(to_unsigned(99, 8)),
			118 => std_logic_vector(to_unsigned(101, 8)),
			119 => std_logic_vector(to_unsigned(129, 8)),
			120 => std_logic_vector(to_unsigned(179, 8)),
			121 => std_logic_vector(to_unsigned(221, 8)),
			122 => std_logic_vector(to_unsigned(224, 8)),
			123 => std_logic_vector(to_unsigned(136, 8)),
			124 => std_logic_vector(to_unsigned(93, 8)),
			125 => std_logic_vector(to_unsigned(124, 8)),
			126 => std_logic_vector(to_unsigned(71, 8)),
			127 => std_logic_vector(to_unsigned(137, 8)),
			128 => std_logic_vector(to_unsigned(227, 8)),
			129 => std_logic_vector(to_unsigned(174, 8)),
			130 => std_logic_vector(to_unsigned(125, 8)),
			131 => std_logic_vector(to_unsigned(115, 8)),
			132 => std_logic_vector(to_unsigned(219, 8)),
			133 => std_logic_vector(to_unsigned(44, 8)),
			134 => std_logic_vector(to_unsigned(242, 8)),
			135 => std_logic_vector(to_unsigned(78, 8)),
			136 => std_logic_vector(to_unsigned(84, 8)),
			137 => std_logic_vector(to_unsigned(219, 8)),
			138 => std_logic_vector(to_unsigned(201, 8)),
			139 => std_logic_vector(to_unsigned(50, 8)),
			140 => std_logic_vector(to_unsigned(249, 8)),
			141 => std_logic_vector(to_unsigned(226, 8)),
			142 => std_logic_vector(to_unsigned(100, 8)),
			143 => std_logic_vector(to_unsigned(69, 8)),
			144 => std_logic_vector(to_unsigned(14, 8)),
			145 => std_logic_vector(to_unsigned(89, 8)),
			146 => std_logic_vector(to_unsigned(46, 8)),
			147 => std_logic_vector(to_unsigned(248, 8)),
			148 => std_logic_vector(to_unsigned(208, 8)),
			149 => std_logic_vector(to_unsigned(125, 8)),
			150 => std_logic_vector(to_unsigned(222, 8)),
			151 => std_logic_vector(to_unsigned(76, 8)),
			152 => std_logic_vector(to_unsigned(128, 8)),
			153 => std_logic_vector(to_unsigned(96, 8)),
			154 => std_logic_vector(to_unsigned(60, 8)),
			155 => std_logic_vector(to_unsigned(226, 8)),
			156 => std_logic_vector(to_unsigned(32, 8)),
			157 => std_logic_vector(to_unsigned(8, 8)),
			158 => std_logic_vector(to_unsigned(13, 8)),
			159 => std_logic_vector(to_unsigned(166, 8)),
			160 => std_logic_vector(to_unsigned(189, 8)),
			161 => std_logic_vector(to_unsigned(101, 8)),
			162 => std_logic_vector(to_unsigned(80, 8)),
			163 => std_logic_vector(to_unsigned(58, 8)),
			164 => std_logic_vector(to_unsigned(1, 8)),
			165 => std_logic_vector(to_unsigned(230, 8)),
			166 => std_logic_vector(to_unsigned(108, 8)),
			167 => std_logic_vector(to_unsigned(40, 8)),
			168 => std_logic_vector(to_unsigned(78, 8)),
			169 => std_logic_vector(to_unsigned(143, 8)),
			170 => std_logic_vector(to_unsigned(9, 8)),
			171 => std_logic_vector(to_unsigned(119, 8)),
			172 => std_logic_vector(to_unsigned(114, 8)),
			173 => std_logic_vector(to_unsigned(163, 8)),
			174 => std_logic_vector(to_unsigned(133, 8)),
			175 => std_logic_vector(to_unsigned(124, 8)),
			176 => std_logic_vector(to_unsigned(190, 8)),
			177 => std_logic_vector(to_unsigned(118, 8)),
			178 => std_logic_vector(to_unsigned(40, 8)),
			179 => std_logic_vector(to_unsigned(53, 8)),
			180 => std_logic_vector(to_unsigned(178, 8)),
			181 => std_logic_vector(to_unsigned(200, 8)),
			182 => std_logic_vector(to_unsigned(29, 8)),
			183 => std_logic_vector(to_unsigned(67, 8)),
			184 => std_logic_vector(to_unsigned(171, 8)),
			185 => std_logic_vector(to_unsigned(71, 8)),
			186 => std_logic_vector(to_unsigned(99, 8)),
			187 => std_logic_vector(to_unsigned(129, 8)),
			188 => std_logic_vector(to_unsigned(110, 8)),
			189 => std_logic_vector(to_unsigned(56, 8)),
			190 => std_logic_vector(to_unsigned(59, 8)),
			191 => std_logic_vector(to_unsigned(36, 8)),
			192 => std_logic_vector(to_unsigned(10, 8)),
			193 => std_logic_vector(to_unsigned(152, 8)),
			194 => std_logic_vector(to_unsigned(6, 8)),
			195 => std_logic_vector(to_unsigned(105, 8)),
			196 => std_logic_vector(to_unsigned(177, 8)),
			197 => std_logic_vector(to_unsigned(56, 8)),
			198 => std_logic_vector(to_unsigned(125, 8)),
			199 => std_logic_vector(to_unsigned(197, 8)),
			200 => std_logic_vector(to_unsigned(228, 8)),
			201 => std_logic_vector(to_unsigned(205, 8)),
			202 => std_logic_vector(to_unsigned(186, 8)),
			203 => std_logic_vector(to_unsigned(84, 8)),
			204 => std_logic_vector(to_unsigned(174, 8)),
			205 => std_logic_vector(to_unsigned(158, 8)),
			206 => std_logic_vector(to_unsigned(41, 8)),
			207 => std_logic_vector(to_unsigned(36, 8)),
			208 => std_logic_vector(to_unsigned(53, 8)),
			209 => std_logic_vector(to_unsigned(97, 8)),
			210 => std_logic_vector(to_unsigned(149, 8)),
			211 => std_logic_vector(to_unsigned(10, 8)),
			212 => std_logic_vector(to_unsigned(116, 8)),
			213 => std_logic_vector(to_unsigned(31, 8)),
			214 => std_logic_vector(to_unsigned(143, 8)),
			215 => std_logic_vector(to_unsigned(145, 8)),
			216 => std_logic_vector(to_unsigned(61, 8)),
			217 => std_logic_vector(to_unsigned(191, 8)),
			218 => std_logic_vector(to_unsigned(143, 8)),
			219 => std_logic_vector(to_unsigned(115, 8)),
			220 => std_logic_vector(to_unsigned(103, 8)),
			221 => std_logic_vector(to_unsigned(228, 8)),
			222 => std_logic_vector(to_unsigned(221, 8)),
			223 => std_logic_vector(to_unsigned(112, 8)),
			224 => std_logic_vector(to_unsigned(172, 8)),
			225 => std_logic_vector(to_unsigned(188, 8)),
			226 => std_logic_vector(to_unsigned(248, 8)),
			227 => std_logic_vector(to_unsigned(174, 8)),
			228 => std_logic_vector(to_unsigned(110, 8)),
			229 => std_logic_vector(to_unsigned(54, 8)),
			230 => std_logic_vector(to_unsigned(53, 8)),
			231 => std_logic_vector(to_unsigned(240, 8)),
			232 => std_logic_vector(to_unsigned(245, 8)),
			233 => std_logic_vector(to_unsigned(188, 8)),
			234 => std_logic_vector(to_unsigned(87, 8)),
			235 => std_logic_vector(to_unsigned(214, 8)),
			236 => std_logic_vector(to_unsigned(20, 8)),
			237 => std_logic_vector(to_unsigned(188, 8)),
			238 => std_logic_vector(to_unsigned(176, 8)),
			239 => std_logic_vector(to_unsigned(187, 8)),
			240 => std_logic_vector(to_unsigned(109, 8)),
			241 => std_logic_vector(to_unsigned(38, 8)),
			242 => std_logic_vector(to_unsigned(247, 8)),
			243 => std_logic_vector(to_unsigned(45, 8)),
			244 => std_logic_vector(to_unsigned(169, 8)),
			245 => std_logic_vector(to_unsigned(114, 8)),
			246 => std_logic_vector(to_unsigned(107, 8)),
			247 => std_logic_vector(to_unsigned(243, 8)),
			248 => std_logic_vector(to_unsigned(157, 8)),
			249 => std_logic_vector(to_unsigned(5, 8)),
			250 => std_logic_vector(to_unsigned(254, 8)),
			251 => std_logic_vector(to_unsigned(130, 8)),
			252 => std_logic_vector(to_unsigned(229, 8)),
			253 => std_logic_vector(to_unsigned(211, 8)),
			254 => std_logic_vector(to_unsigned(89, 8)),
			255 => std_logic_vector(to_unsigned(157, 8)),
			256 => std_logic_vector(to_unsigned(6, 8)),
			257 => std_logic_vector(to_unsigned(237, 8)),
			258 => std_logic_vector(to_unsigned(61, 8)),
			259 => std_logic_vector(to_unsigned(252, 8)),
			260 => std_logic_vector(to_unsigned(5, 8)),
			261 => std_logic_vector(to_unsigned(174, 8)),
			262 => std_logic_vector(to_unsigned(30, 8)),
			263 => std_logic_vector(to_unsigned(200, 8)),
			264 => std_logic_vector(to_unsigned(19, 8)),
			265 => std_logic_vector(to_unsigned(137, 8)),
			266 => std_logic_vector(to_unsigned(108, 8)),
			267 => std_logic_vector(to_unsigned(89, 8)),
			268 => std_logic_vector(to_unsigned(183, 8)),
			269 => std_logic_vector(to_unsigned(106, 8)),
			270 => std_logic_vector(to_unsigned(176, 8)),
			271 => std_logic_vector(to_unsigned(245, 8)),
			272 => std_logic_vector(to_unsigned(114, 8)),
			273 => std_logic_vector(to_unsigned(151, 8)),
			274 => std_logic_vector(to_unsigned(29, 8)),
			275 => std_logic_vector(to_unsigned(189, 8)),
			276 => std_logic_vector(to_unsigned(134, 8)),
			277 => std_logic_vector(to_unsigned(158, 8)),
			278 => std_logic_vector(to_unsigned(89, 8)),
			279 => std_logic_vector(to_unsigned(142, 8)),
			280 => std_logic_vector(to_unsigned(206, 8)),
			281 => std_logic_vector(to_unsigned(190, 8)),
			282 => std_logic_vector(to_unsigned(89, 8)),
			283 => std_logic_vector(to_unsigned(5, 8)),
			284 => std_logic_vector(to_unsigned(191, 8)),
			285 => std_logic_vector(to_unsigned(46, 8)),
			286 => std_logic_vector(to_unsigned(154, 8)),
			287 => std_logic_vector(to_unsigned(109, 8)),
			288 => std_logic_vector(to_unsigned(67, 8)),
			289 => std_logic_vector(to_unsigned(237, 8)),
			290 => std_logic_vector(to_unsigned(139, 8)),
			291 => std_logic_vector(to_unsigned(201, 8)),
			292 => std_logic_vector(to_unsigned(195, 8)),
			293 => std_logic_vector(to_unsigned(147, 8)),
			294 => std_logic_vector(to_unsigned(67, 8)),
			295 => std_logic_vector(to_unsigned(214, 8)),
			296 => std_logic_vector(to_unsigned(209, 8)),
			297 => std_logic_vector(to_unsigned(230, 8)),
			298 => std_logic_vector(to_unsigned(80, 8)),
			299 => std_logic_vector(to_unsigned(25, 8)),
			300 => std_logic_vector(to_unsigned(179, 8)),
			301 => std_logic_vector(to_unsigned(113, 8)),
			302 => std_logic_vector(to_unsigned(13, 8)),
			303 => std_logic_vector(to_unsigned(205, 8)),
			304 => std_logic_vector(to_unsigned(52, 8)),
			305 => std_logic_vector(to_unsigned(177, 8)),
			306 => std_logic_vector(to_unsigned(169, 8)),
			307 => std_logic_vector(to_unsigned(157, 8)),
			308 => std_logic_vector(to_unsigned(246, 8)),
			309 => std_logic_vector(to_unsigned(210, 8)),
			310 => std_logic_vector(to_unsigned(128, 8)),
			311 => std_logic_vector(to_unsigned(36, 8)),
			312 => std_logic_vector(to_unsigned(130, 8)),
			313 => std_logic_vector(to_unsigned(86, 8)),
			314 => std_logic_vector(to_unsigned(162, 8)),
			315 => std_logic_vector(to_unsigned(106, 8)),
			316 => std_logic_vector(to_unsigned(165, 8)),
			317 => std_logic_vector(to_unsigned(149, 8)),
			318 => std_logic_vector(to_unsigned(93, 8)),
			319 => std_logic_vector(to_unsigned(145, 8)),
			320 => std_logic_vector(to_unsigned(139, 8)),
			321 => std_logic_vector(to_unsigned(0, 8)),
			322 => std_logic_vector(to_unsigned(238, 8)),
			323 => std_logic_vector(to_unsigned(78, 8)),
			324 => std_logic_vector(to_unsigned(28, 8)),
			325 => std_logic_vector(to_unsigned(193, 8)),
			326 => std_logic_vector(to_unsigned(134, 8)),
			327 => std_logic_vector(to_unsigned(227, 8)),
			328 => std_logic_vector(to_unsigned(121, 8)),
			329 => std_logic_vector(to_unsigned(111, 8)),
			330 => std_logic_vector(to_unsigned(252, 8)),
			331 => std_logic_vector(to_unsigned(149, 8)),
			332 => std_logic_vector(to_unsigned(3, 8)),
			333 => std_logic_vector(to_unsigned(182, 8)),
			334 => std_logic_vector(to_unsigned(206, 8)),
			335 => std_logic_vector(to_unsigned(14, 8)),
			336 => std_logic_vector(to_unsigned(15, 8)),
			337 => std_logic_vector(to_unsigned(210, 8)),
			338 => std_logic_vector(to_unsigned(90, 8)),
			339 => std_logic_vector(to_unsigned(253, 8)),
			340 => std_logic_vector(to_unsigned(31, 8)),
			341 => std_logic_vector(to_unsigned(14, 8)),
			342 => std_logic_vector(to_unsigned(119, 8)),
			343 => std_logic_vector(to_unsigned(35, 8)),
			344 => std_logic_vector(to_unsigned(119, 8)),
			345 => std_logic_vector(to_unsigned(239, 8)),
			346 => std_logic_vector(to_unsigned(69, 8)),
			347 => std_logic_vector(to_unsigned(81, 8)),
			348 => std_logic_vector(to_unsigned(248, 8)),
			349 => std_logic_vector(to_unsigned(238, 8)),
			350 => std_logic_vector(to_unsigned(183, 8)),
			351 => std_logic_vector(to_unsigned(34, 8)),
			352 => std_logic_vector(to_unsigned(116, 8)),
			353 => std_logic_vector(to_unsigned(49, 8)),
			354 => std_logic_vector(to_unsigned(38, 8)),
			355 => std_logic_vector(to_unsigned(45, 8)),
			356 => std_logic_vector(to_unsigned(221, 8)),
			357 => std_logic_vector(to_unsigned(184, 8)),
			358 => std_logic_vector(to_unsigned(172, 8)),
			359 => std_logic_vector(to_unsigned(212, 8)),
			360 => std_logic_vector(to_unsigned(206, 8)),
			361 => std_logic_vector(to_unsigned(189, 8)),
			362 => std_logic_vector(to_unsigned(44, 8)),
			363 => std_logic_vector(to_unsigned(255, 8)),
			364 => std_logic_vector(to_unsigned(252, 8)),
			365 => std_logic_vector(to_unsigned(72, 8)),
			366 => std_logic_vector(to_unsigned(187, 8)),
			367 => std_logic_vector(to_unsigned(231, 8)),
			368 => std_logic_vector(to_unsigned(191, 8)),
			369 => std_logic_vector(to_unsigned(156, 8)),
			370 => std_logic_vector(to_unsigned(237, 8)),
			371 => std_logic_vector(to_unsigned(204, 8)),
			372 => std_logic_vector(to_unsigned(241, 8)),
			373 => std_logic_vector(to_unsigned(214, 8)),
			374 => std_logic_vector(to_unsigned(117, 8)),
			375 => std_logic_vector(to_unsigned(120, 8)),
			376 => std_logic_vector(to_unsigned(172, 8)),
			377 => std_logic_vector(to_unsigned(119, 8)),
			378 => std_logic_vector(to_unsigned(193, 8)),
			379 => std_logic_vector(to_unsigned(50, 8)),
			380 => std_logic_vector(to_unsigned(68, 8)),
			381 => std_logic_vector(to_unsigned(99, 8)),
			382 => std_logic_vector(to_unsigned(160, 8)),
			383 => std_logic_vector(to_unsigned(192, 8)),
			384 => std_logic_vector(to_unsigned(146, 8)),
			385 => std_logic_vector(to_unsigned(213, 8)),
			386 => std_logic_vector(to_unsigned(159, 8)),
			387 => std_logic_vector(to_unsigned(196, 8)),
			388 => std_logic_vector(to_unsigned(56, 8)),
			389 => std_logic_vector(to_unsigned(192, 8)),
			390 => std_logic_vector(to_unsigned(220, 8)),
			391 => std_logic_vector(to_unsigned(69, 8)),
			392 => std_logic_vector(to_unsigned(135, 8)),
			393 => std_logic_vector(to_unsigned(168, 8)),
			394 => std_logic_vector(to_unsigned(32, 8)),
			395 => std_logic_vector(to_unsigned(50, 8)),
			396 => std_logic_vector(to_unsigned(74, 8)),
			397 => std_logic_vector(to_unsigned(74, 8)),
			398 => std_logic_vector(to_unsigned(179, 8)),
			399 => std_logic_vector(to_unsigned(119, 8)),
			400 => std_logic_vector(to_unsigned(76, 8)),
			401 => std_logic_vector(to_unsigned(217, 8)),
			402 => std_logic_vector(to_unsigned(185, 8)),
			403 => std_logic_vector(to_unsigned(108, 8)),
			404 => std_logic_vector(to_unsigned(238, 8)),
			405 => std_logic_vector(to_unsigned(53, 8)),
			406 => std_logic_vector(to_unsigned(216, 8)),
			407 => std_logic_vector(to_unsigned(123, 8)),
			408 => std_logic_vector(to_unsigned(97, 8)),
			409 => std_logic_vector(to_unsigned(30, 8)),
			410 => std_logic_vector(to_unsigned(106, 8)),
			411 => std_logic_vector(to_unsigned(222, 8)),
			412 => std_logic_vector(to_unsigned(172, 8)),
			413 => std_logic_vector(to_unsigned(64, 8)),
			414 => std_logic_vector(to_unsigned(139, 8)),
			415 => std_logic_vector(to_unsigned(90, 8)),
			416 => std_logic_vector(to_unsigned(222, 8)),
			417 => std_logic_vector(to_unsigned(156, 8)),
			418 => std_logic_vector(to_unsigned(228, 8)),
			419 => std_logic_vector(to_unsigned(61, 8)),
			420 => std_logic_vector(to_unsigned(81, 8)),
			421 => std_logic_vector(to_unsigned(203, 8)),
			422 => std_logic_vector(to_unsigned(20, 8)),
			423 => std_logic_vector(to_unsigned(179, 8)),
			424 => std_logic_vector(to_unsigned(86, 8)),
			425 => std_logic_vector(to_unsigned(208, 8)),
			426 => std_logic_vector(to_unsigned(52, 8)),
			427 => std_logic_vector(to_unsigned(228, 8)),
			428 => std_logic_vector(to_unsigned(127, 8)),
			429 => std_logic_vector(to_unsigned(60, 8)),
			430 => std_logic_vector(to_unsigned(119, 8)),
			431 => std_logic_vector(to_unsigned(196, 8)),
			432 => std_logic_vector(to_unsigned(55, 8)),
			433 => std_logic_vector(to_unsigned(206, 8)),
			434 => std_logic_vector(to_unsigned(57, 8)),
			435 => std_logic_vector(to_unsigned(114, 8)),
			436 => std_logic_vector(to_unsigned(21, 8)),
			437 => std_logic_vector(to_unsigned(216, 8)),
			438 => std_logic_vector(to_unsigned(133, 8)),
			439 => std_logic_vector(to_unsigned(28, 8)),
			440 => std_logic_vector(to_unsigned(68, 8)),
			441 => std_logic_vector(to_unsigned(120, 8)),
			442 => std_logic_vector(to_unsigned(238, 8)),
			443 => std_logic_vector(to_unsigned(204, 8)),
			444 => std_logic_vector(to_unsigned(190, 8)),
			445 => std_logic_vector(to_unsigned(208, 8)),
			446 => std_logic_vector(to_unsigned(51, 8)),
			447 => std_logic_vector(to_unsigned(87, 8)),
			448 => std_logic_vector(to_unsigned(232, 8)),
			449 => std_logic_vector(to_unsigned(209, 8)),
			450 => std_logic_vector(to_unsigned(52, 8)),
			451 => std_logic_vector(to_unsigned(2, 8)),
			452 => std_logic_vector(to_unsigned(203, 8)),
			453 => std_logic_vector(to_unsigned(81, 8)),
			454 => std_logic_vector(to_unsigned(3, 8)),
			455 => std_logic_vector(to_unsigned(226, 8)),
			456 => std_logic_vector(to_unsigned(227, 8)),
			457 => std_logic_vector(to_unsigned(139, 8)),
			458 => std_logic_vector(to_unsigned(114, 8)),
			459 => std_logic_vector(to_unsigned(33, 8)),
			460 => std_logic_vector(to_unsigned(169, 8)),
			461 => std_logic_vector(to_unsigned(207, 8)),
			462 => std_logic_vector(to_unsigned(172, 8)),
			463 => std_logic_vector(to_unsigned(79, 8)),
			464 => std_logic_vector(to_unsigned(251, 8)),
			465 => std_logic_vector(to_unsigned(36, 8)),
			466 => std_logic_vector(to_unsigned(225, 8)),
			467 => std_logic_vector(to_unsigned(206, 8)),
			468 => std_logic_vector(to_unsigned(68, 8)),
			469 => std_logic_vector(to_unsigned(237, 8)),
			470 => std_logic_vector(to_unsigned(233, 8)),
			471 => std_logic_vector(to_unsigned(204, 8)),
			472 => std_logic_vector(to_unsigned(172, 8)),
			473 => std_logic_vector(to_unsigned(159, 8)),
			474 => std_logic_vector(to_unsigned(98, 8)),
			475 => std_logic_vector(to_unsigned(39, 8)),
			476 => std_logic_vector(to_unsigned(216, 8)),
			477 => std_logic_vector(to_unsigned(83, 8)),
			478 => std_logic_vector(to_unsigned(240, 8)),
			479 => std_logic_vector(to_unsigned(232, 8)),
			480 => std_logic_vector(to_unsigned(241, 8)),
			481 => std_logic_vector(to_unsigned(208, 8)),
			482 => std_logic_vector(to_unsigned(59, 8)),
			483 => std_logic_vector(to_unsigned(1, 8)),
			484 => std_logic_vector(to_unsigned(22, 8)),
			485 => std_logic_vector(to_unsigned(157, 8)),
			486 => std_logic_vector(to_unsigned(108, 8)),
			487 => std_logic_vector(to_unsigned(82, 8)),
			488 => std_logic_vector(to_unsigned(254, 8)),
			489 => std_logic_vector(to_unsigned(207, 8)),
			490 => std_logic_vector(to_unsigned(99, 8)),
			491 => std_logic_vector(to_unsigned(144, 8)),
			492 => std_logic_vector(to_unsigned(211, 8)),
			493 => std_logic_vector(to_unsigned(77, 8)),
			494 => std_logic_vector(to_unsigned(186, 8)),
			495 => std_logic_vector(to_unsigned(128, 8)),
			496 => std_logic_vector(to_unsigned(243, 8)),
			497 => std_logic_vector(to_unsigned(59, 8)),
			498 => std_logic_vector(to_unsigned(13, 8)),
			499 => std_logic_vector(to_unsigned(108, 8)),
			500 => std_logic_vector(to_unsigned(151, 8)),
			501 => std_logic_vector(to_unsigned(51, 8)),
			502 => std_logic_vector(to_unsigned(75, 8)),
			503 => std_logic_vector(to_unsigned(71, 8)),
			504 => std_logic_vector(to_unsigned(98, 8)),
			505 => std_logic_vector(to_unsigned(160, 8)),
			506 => std_logic_vector(to_unsigned(214, 8)),
			507 => std_logic_vector(to_unsigned(161, 8)),
			508 => std_logic_vector(to_unsigned(221, 8)),
			509 => std_logic_vector(to_unsigned(104, 8)),
			510 => std_logic_vector(to_unsigned(128, 8)),
			511 => std_logic_vector(to_unsigned(126, 8)),
			512 => std_logic_vector(to_unsigned(10, 8)),
			513 => std_logic_vector(to_unsigned(219, 8)),
			514 => std_logic_vector(to_unsigned(96, 8)),
			515 => std_logic_vector(to_unsigned(96, 8)),
			516 => std_logic_vector(to_unsigned(230, 8)),
			517 => std_logic_vector(to_unsigned(91, 8)),
			518 => std_logic_vector(to_unsigned(35, 8)),
			519 => std_logic_vector(to_unsigned(217, 8)),
			520 => std_logic_vector(to_unsigned(161, 8)),
			521 => std_logic_vector(to_unsigned(238, 8)),
			522 => std_logic_vector(to_unsigned(238, 8)),
			523 => std_logic_vector(to_unsigned(71, 8)),
			524 => std_logic_vector(to_unsigned(59, 8)),
			525 => std_logic_vector(to_unsigned(163, 8)),
			526 => std_logic_vector(to_unsigned(193, 8)),
			527 => std_logic_vector(to_unsigned(146, 8)),
			528 => std_logic_vector(to_unsigned(1, 8)),
			529 => std_logic_vector(to_unsigned(30, 8)),
			530 => std_logic_vector(to_unsigned(232, 8)),
			531 => std_logic_vector(to_unsigned(239, 8)),
			532 => std_logic_vector(to_unsigned(222, 8)),
			533 => std_logic_vector(to_unsigned(122, 8)),
			534 => std_logic_vector(to_unsigned(177, 8)),
			535 => std_logic_vector(to_unsigned(0, 8)),
			536 => std_logic_vector(to_unsigned(186, 8)),
			537 => std_logic_vector(to_unsigned(18, 8)),
			538 => std_logic_vector(to_unsigned(213, 8)),
			539 => std_logic_vector(to_unsigned(219, 8)),
			540 => std_logic_vector(to_unsigned(69, 8)),
			541 => std_logic_vector(to_unsigned(134, 8)),
			542 => std_logic_vector(to_unsigned(177, 8)),
			543 => std_logic_vector(to_unsigned(233, 8)),
			544 => std_logic_vector(to_unsigned(188, 8)),
			545 => std_logic_vector(to_unsigned(174, 8)),
			546 => std_logic_vector(to_unsigned(139, 8)),
			547 => std_logic_vector(to_unsigned(164, 8)),
			548 => std_logic_vector(to_unsigned(59, 8)),
			549 => std_logic_vector(to_unsigned(203, 8)),
			550 => std_logic_vector(to_unsigned(195, 8)),
			551 => std_logic_vector(to_unsigned(192, 8)),
			552 => std_logic_vector(to_unsigned(17, 8)),
			553 => std_logic_vector(to_unsigned(142, 8)),
			554 => std_logic_vector(to_unsigned(60, 8)),
			555 => std_logic_vector(to_unsigned(242, 8)),
			556 => std_logic_vector(to_unsigned(237, 8)),
			557 => std_logic_vector(to_unsigned(252, 8)),
			558 => std_logic_vector(to_unsigned(143, 8)),
			559 => std_logic_vector(to_unsigned(106, 8)),
			560 => std_logic_vector(to_unsigned(161, 8)),
			561 => std_logic_vector(to_unsigned(153, 8)),
			562 => std_logic_vector(to_unsigned(5, 8)),
			563 => std_logic_vector(to_unsigned(133, 8)),
			564 => std_logic_vector(to_unsigned(154, 8)),
			565 => std_logic_vector(to_unsigned(210, 8)),
			566 => std_logic_vector(to_unsigned(204, 8)),
			567 => std_logic_vector(to_unsigned(105, 8)),
			568 => std_logic_vector(to_unsigned(86, 8)),
			569 => std_logic_vector(to_unsigned(243, 8)),
			570 => std_logic_vector(to_unsigned(106, 8)),
			571 => std_logic_vector(to_unsigned(2, 8)),
			572 => std_logic_vector(to_unsigned(5, 8)),
			573 => std_logic_vector(to_unsigned(230, 8)),
			574 => std_logic_vector(to_unsigned(65, 8)),
			575 => std_logic_vector(to_unsigned(202, 8)),
			576 => std_logic_vector(to_unsigned(252, 8)),
			577 => std_logic_vector(to_unsigned(137, 8)),
			578 => std_logic_vector(to_unsigned(13, 8)),
			579 => std_logic_vector(to_unsigned(227, 8)),
			580 => std_logic_vector(to_unsigned(75, 8)),
			581 => std_logic_vector(to_unsigned(69, 8)),
			582 => std_logic_vector(to_unsigned(202, 8)),
			583 => std_logic_vector(to_unsigned(31, 8)),
			584 => std_logic_vector(to_unsigned(63, 8)),
			585 => std_logic_vector(to_unsigned(140, 8)),
			586 => std_logic_vector(to_unsigned(65, 8)),
			587 => std_logic_vector(to_unsigned(247, 8)),
			588 => std_logic_vector(to_unsigned(162, 8)),
			589 => std_logic_vector(to_unsigned(7, 8)),
			590 => std_logic_vector(to_unsigned(74, 8)),
			591 => std_logic_vector(to_unsigned(105, 8)),
			592 => std_logic_vector(to_unsigned(8, 8)),
			593 => std_logic_vector(to_unsigned(190, 8)),
			594 => std_logic_vector(to_unsigned(75, 8)),
			595 => std_logic_vector(to_unsigned(52, 8)),
			596 => std_logic_vector(to_unsigned(169, 8)),
			597 => std_logic_vector(to_unsigned(183, 8)),
			598 => std_logic_vector(to_unsigned(54, 8)),
			599 => std_logic_vector(to_unsigned(252, 8)),
			600 => std_logic_vector(to_unsigned(37, 8)),
			601 => std_logic_vector(to_unsigned(228, 8)),
			602 => std_logic_vector(to_unsigned(207, 8)),
			603 => std_logic_vector(to_unsigned(200, 8)),
			604 => std_logic_vector(to_unsigned(98, 8)),
			605 => std_logic_vector(to_unsigned(32, 8)),
			606 => std_logic_vector(to_unsigned(150, 8)),
			607 => std_logic_vector(to_unsigned(101, 8)),
			608 => std_logic_vector(to_unsigned(77, 8)),
			609 => std_logic_vector(to_unsigned(136, 8)),
			610 => std_logic_vector(to_unsigned(129, 8)),
			611 => std_logic_vector(to_unsigned(151, 8)),
			612 => std_logic_vector(to_unsigned(22, 8)),
			613 => std_logic_vector(to_unsigned(208, 8)),
			614 => std_logic_vector(to_unsigned(206, 8)),
			615 => std_logic_vector(to_unsigned(20, 8)),
			616 => std_logic_vector(to_unsigned(160, 8)),
			617 => std_logic_vector(to_unsigned(10, 8)),
			618 => std_logic_vector(to_unsigned(204, 8)),
			619 => std_logic_vector(to_unsigned(4, 8)),
			620 => std_logic_vector(to_unsigned(36, 8)),
			621 => std_logic_vector(to_unsigned(146, 8)),
			622 => std_logic_vector(to_unsigned(65, 8)),
			623 => std_logic_vector(to_unsigned(24, 8)),
			624 => std_logic_vector(to_unsigned(29, 8)),
			625 => std_logic_vector(to_unsigned(201, 8)),
			626 => std_logic_vector(to_unsigned(247, 8)),
			627 => std_logic_vector(to_unsigned(254, 8)),
			628 => std_logic_vector(to_unsigned(219, 8)),
			629 => std_logic_vector(to_unsigned(220, 8)),
			630 => std_logic_vector(to_unsigned(56, 8)),
			631 => std_logic_vector(to_unsigned(3, 8)),
			632 => std_logic_vector(to_unsigned(233, 8)),
			633 => std_logic_vector(to_unsigned(65, 8)),
			634 => std_logic_vector(to_unsigned(211, 8)),
			635 => std_logic_vector(to_unsigned(231, 8)),
			636 => std_logic_vector(to_unsigned(18, 8)),
			637 => std_logic_vector(to_unsigned(0, 8)),
			638 => std_logic_vector(to_unsigned(135, 8)),
			639 => std_logic_vector(to_unsigned(20, 8)),
			others => (others => '0'));                       

component project_reti_logiche is
port (
      i_clk         : in  std_logic;
      i_rst         : in  std_logic;
      i_start       : in  std_logic;
      i_data        : in  std_logic_vector(7 downto 0);
      o_address     : out std_logic_vector(15 downto 0);
      o_done        : out std_logic;
      o_en          : out std_logic;
      o_we          : out std_logic;
      o_data        : out std_logic_vector (7 downto 0)
      );
end component project_reti_logiche;


begin
UUT: project_reti_logiche
port map (
          i_clk      	=> tb_clk,
          i_rst      	=> tb_rst,
          i_start       => tb_start,
          i_data    	=> mem_o_data,
          o_address  	=> mem_address,
          o_done      	=> tb_done,
          o_en   	=> enable_wire,
          o_we 		=> mem_we,
          o_data    	=> mem_i_data
          );

p_CLK_GEN : process is
begin
    wait for c_CLOCK_PERIOD/2;
    tb_clk <= not tb_clk;
end process p_CLK_GEN;


MEM : process(tb_clk)
begin
    if tb_clk'event and tb_clk = '1' then
        if enable_wire = '1' then
            if mem_we = '1' then
                RAM(conv_integer(mem_address))  <= mem_i_data;
                mem_o_data                      <= mem_i_data after 1 ns;
            else
                mem_o_data <= RAM(conv_integer(mem_address)) after 1 ns;
            end if;
        end if;
    end if;
end process;


test : process is
begin 
    wait for 100 ns;
    wait for c_CLOCK_PERIOD;
    tb_rst <= '1';
    wait for c_CLOCK_PERIOD;
    wait for 100 ns;
    tb_rst <= '0';
    wait for c_CLOCK_PERIOD;
    wait for 100 ns;
    tb_start <= '1';
    wait for c_CLOCK_PERIOD;
    wait until tb_done = '1';
    wait for c_CLOCK_PERIOD;
    tb_start <= '0';
    wait until tb_done = '0';
    wait for 100 ns;
    
    assert RAM(640) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(640))))  severity failure;
	assert RAM(641) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(641))))  severity failure;
	assert RAM(642) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(642))))  severity failure;
	assert RAM(643) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(643))))  severity failure;
	assert RAM(644) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(644))))  severity failure;
	assert RAM(645) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(645))))  severity failure;
	assert RAM(646) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(646))))  severity failure;
	assert RAM(647) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(647))))  severity failure;
	assert RAM(648) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(648))))  severity failure;
	assert RAM(649) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(649))))  severity failure;
	assert RAM(650) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(650))))  severity failure;
	assert RAM(651) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(651))))  severity failure;
	assert RAM(652) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(652))))  severity failure;
	assert RAM(653) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(653))))  severity failure;
	assert RAM(654) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(654))))  severity failure;
	assert RAM(655) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(655))))  severity failure;
	assert RAM(656) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(656))))  severity failure;
	assert RAM(657) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(657))))  severity failure;
	assert RAM(658) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(658))))  severity failure;
	assert RAM(659) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(659))))  severity failure;
	assert RAM(660) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(660))))  severity failure;
	assert RAM(661) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(661))))  severity failure;
	assert RAM(662) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(662))))  severity failure;
	assert RAM(663) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(663))))  severity failure;
	assert RAM(664) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(664))))  severity failure;
	assert RAM(665) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(665))))  severity failure;
	assert RAM(666) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(666))))  severity failure;
	assert RAM(667) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(667))))  severity failure;
	assert RAM(668) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(668))))  severity failure;
	assert RAM(669) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(669))))  severity failure;
	assert RAM(670) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(670))))  severity failure;
	assert RAM(671) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(671))))  severity failure;
	assert RAM(672) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(672))))  severity failure;
	assert RAM(673) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(673))))  severity failure;
	assert RAM(674) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(674))))  severity failure;
	assert RAM(675) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(675))))  severity failure;
	assert RAM(676) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(676))))  severity failure;
	assert RAM(677) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(677))))  severity failure;
	assert RAM(678) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(678))))  severity failure;
	assert RAM(679) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(679))))  severity failure;
	assert RAM(680) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(680))))  severity failure;
	assert RAM(681) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(681))))  severity failure;
	assert RAM(682) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(682))))  severity failure;
	assert RAM(683) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(683))))  severity failure;
	assert RAM(684) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(684))))  severity failure;
	assert RAM(685) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(685))))  severity failure;
	assert RAM(686) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(686))))  severity failure;
	assert RAM(687) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(687))))  severity failure;
	assert RAM(688) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(688))))  severity failure;
	assert RAM(689) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(689))))  severity failure;
	assert RAM(690) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(690))))  severity failure;
	assert RAM(691) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(691))))  severity failure;
	assert RAM(692) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(692))))  severity failure;
	assert RAM(693) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(693))))  severity failure;
	assert RAM(694) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(694))))  severity failure;
	assert RAM(695) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(695))))  severity failure;
	assert RAM(696) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(696))))  severity failure;
	assert RAM(697) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(697))))  severity failure;
	assert RAM(698) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(698))))  severity failure;
	assert RAM(699) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(699))))  severity failure;
	assert RAM(700) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(700))))  severity failure;
	assert RAM(701) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(701))))  severity failure;
	assert RAM(702) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(702))))  severity failure;
	assert RAM(703) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(703))))  severity failure;
	assert RAM(704) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(704))))  severity failure;
	assert RAM(705) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(705))))  severity failure;
	assert RAM(706) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(706))))  severity failure;
	assert RAM(707) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(707))))  severity failure;
	assert RAM(708) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(708))))  severity failure;
	assert RAM(709) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(709))))  severity failure;
	assert RAM(710) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(710))))  severity failure;
	assert RAM(711) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(711))))  severity failure;
	assert RAM(712) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(712))))  severity failure;
	assert RAM(713) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(713))))  severity failure;
	assert RAM(714) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(714))))  severity failure;
	assert RAM(715) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(715))))  severity failure;
	assert RAM(716) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(716))))  severity failure;
	assert RAM(717) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(717))))  severity failure;
	assert RAM(718) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(718))))  severity failure;
	assert RAM(719) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(719))))  severity failure;
	assert RAM(720) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(720))))  severity failure;
	assert RAM(721) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(721))))  severity failure;
	assert RAM(722) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(722))))  severity failure;
	assert RAM(723) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(723))))  severity failure;
	assert RAM(724) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(724))))  severity failure;
	assert RAM(725) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(725))))  severity failure;
	assert RAM(726) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(726))))  severity failure;
	assert RAM(727) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(727))))  severity failure;
	assert RAM(728) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(728))))  severity failure;
	assert RAM(729) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(729))))  severity failure;
	assert RAM(730) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(730))))  severity failure;
	assert RAM(731) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(731))))  severity failure;
	assert RAM(732) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(732))))  severity failure;
	assert RAM(733) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(733))))  severity failure;
	assert RAM(734) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(734))))  severity failure;
	assert RAM(735) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(735))))  severity failure;
	assert RAM(736) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(736))))  severity failure;
	assert RAM(737) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(737))))  severity failure;
	assert RAM(738) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(738))))  severity failure;
	assert RAM(739) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(739))))  severity failure;
	assert RAM(740) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(740))))  severity failure;
	assert RAM(741) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(741))))  severity failure;
	assert RAM(742) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(742))))  severity failure;
	assert RAM(743) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(743))))  severity failure;
	assert RAM(744) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(744))))  severity failure;
	assert RAM(745) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(745))))  severity failure;
	assert RAM(746) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(746))))  severity failure;
	assert RAM(747) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(747))))  severity failure;
	assert RAM(748) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(748))))  severity failure;
	assert RAM(749) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(749))))  severity failure;
	assert RAM(750) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(750))))  severity failure;
	assert RAM(751) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(751))))  severity failure;
	assert RAM(752) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(752))))  severity failure;
	assert RAM(753) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(753))))  severity failure;
	assert RAM(754) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(754))))  severity failure;
	assert RAM(755) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(755))))  severity failure;
	assert RAM(756) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(756))))  severity failure;
	assert RAM(757) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(757))))  severity failure;
	assert RAM(758) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(758))))  severity failure;
	assert RAM(759) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(759))))  severity failure;
	assert RAM(760) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(760))))  severity failure;
	assert RAM(761) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(761))))  severity failure;
	assert RAM(762) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(762))))  severity failure;
	assert RAM(763) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(763))))  severity failure;
	assert RAM(764) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(764))))  severity failure;
	assert RAM(765) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(765))))  severity failure;
	assert RAM(766) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(766))))  severity failure;
	assert RAM(767) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(767))))  severity failure;
	assert RAM(768) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(768))))  severity failure;
	assert RAM(769) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(769))))  severity failure;
	assert RAM(770) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(770))))  severity failure;
	assert RAM(771) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(771))))  severity failure;
	assert RAM(772) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(772))))  severity failure;
	assert RAM(773) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(773))))  severity failure;
	assert RAM(774) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(774))))  severity failure;
	assert RAM(775) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(775))))  severity failure;
	assert RAM(776) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(776))))  severity failure;
	assert RAM(777) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(777))))  severity failure;
	assert RAM(778) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(778))))  severity failure;
	assert RAM(779) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(779))))  severity failure;
	assert RAM(780) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(780))))  severity failure;
	assert RAM(781) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(781))))  severity failure;
	assert RAM(782) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(782))))  severity failure;
	assert RAM(783) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(783))))  severity failure;
	assert RAM(784) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(784))))  severity failure;
	assert RAM(785) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(785))))  severity failure;
	assert RAM(786) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(786))))  severity failure;
	assert RAM(787) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(787))))  severity failure;
	assert RAM(788) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(788))))  severity failure;
	assert RAM(789) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(789))))  severity failure;
	assert RAM(790) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(790))))  severity failure;
	assert RAM(791) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(791))))  severity failure;
	assert RAM(792) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(792))))  severity failure;
	assert RAM(793) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(793))))  severity failure;
	assert RAM(794) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(794))))  severity failure;
	assert RAM(795) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(795))))  severity failure;
	assert RAM(796) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(796))))  severity failure;
	assert RAM(797) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(797))))  severity failure;
	assert RAM(798) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(798))))  severity failure;
	assert RAM(799) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(799))))  severity failure;
	assert RAM(800) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(800))))  severity failure;
	assert RAM(801) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(801))))  severity failure;
	assert RAM(802) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(802))))  severity failure;
	assert RAM(803) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(803))))  severity failure;
	assert RAM(804) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(804))))  severity failure;
	assert RAM(805) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(805))))  severity failure;
	assert RAM(806) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(806))))  severity failure;
	assert RAM(807) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(807))))  severity failure;
	assert RAM(808) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(808))))  severity failure;
	assert RAM(809) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(809))))  severity failure;
	assert RAM(810) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(810))))  severity failure;
	assert RAM(811) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(811))))  severity failure;
	assert RAM(812) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(812))))  severity failure;
	assert RAM(813) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(813))))  severity failure;
	assert RAM(814) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(814))))  severity failure;
	assert RAM(815) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(815))))  severity failure;
	assert RAM(816) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(816))))  severity failure;
	assert RAM(817) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(817))))  severity failure;
	assert RAM(818) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(818))))  severity failure;
	assert RAM(819) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(819))))  severity failure;
	assert RAM(820) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(820))))  severity failure;
	assert RAM(821) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(821))))  severity failure;
	assert RAM(822) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(822))))  severity failure;
	assert RAM(823) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(823))))  severity failure;
	assert RAM(824) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(824))))  severity failure;
	assert RAM(825) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(825))))  severity failure;
	assert RAM(826) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(826))))  severity failure;
	assert RAM(827) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(827))))  severity failure;
	assert RAM(828) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(828))))  severity failure;
	assert RAM(829) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(829))))  severity failure;
	assert RAM(830) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(830))))  severity failure;
	assert RAM(831) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(831))))  severity failure;
	assert RAM(832) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(832))))  severity failure;
	assert RAM(833) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(833))))  severity failure;
	assert RAM(834) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(834))))  severity failure;
	assert RAM(835) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(835))))  severity failure;
	assert RAM(836) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(836))))  severity failure;
	assert RAM(837) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(837))))  severity failure;
	assert RAM(838) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(838))))  severity failure;
	assert RAM(839) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(839))))  severity failure;
	assert RAM(840) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(840))))  severity failure;
	assert RAM(841) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(841))))  severity failure;
	assert RAM(842) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(842))))  severity failure;
	assert RAM(843) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(843))))  severity failure;
	assert RAM(844) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(844))))  severity failure;
	assert RAM(845) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(845))))  severity failure;
	assert RAM(846) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(846))))  severity failure;
	assert RAM(847) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(847))))  severity failure;
	assert RAM(848) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(848))))  severity failure;
	assert RAM(849) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(849))))  severity failure;
	assert RAM(850) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(850))))  severity failure;
	assert RAM(851) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(851))))  severity failure;
	assert RAM(852) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(852))))  severity failure;
	assert RAM(853) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(853))))  severity failure;
	assert RAM(854) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(854))))  severity failure;
	assert RAM(855) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(855))))  severity failure;
	assert RAM(856) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(856))))  severity failure;
	assert RAM(857) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(857))))  severity failure;
	assert RAM(858) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(858))))  severity failure;
	assert RAM(859) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(859))))  severity failure;
	assert RAM(860) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(860))))  severity failure;
	assert RAM(861) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(861))))  severity failure;
	assert RAM(862) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(862))))  severity failure;
	assert RAM(863) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(863))))  severity failure;
	assert RAM(864) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(864))))  severity failure;
	assert RAM(865) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(865))))  severity failure;
	assert RAM(866) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(866))))  severity failure;
	assert RAM(867) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(867))))  severity failure;
	assert RAM(868) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(868))))  severity failure;
	assert RAM(869) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(869))))  severity failure;
	assert RAM(870) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(870))))  severity failure;
	assert RAM(871) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(871))))  severity failure;
	assert RAM(872) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(872))))  severity failure;
	assert RAM(873) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(873))))  severity failure;
	assert RAM(874) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(874))))  severity failure;
	assert RAM(875) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(875))))  severity failure;
	assert RAM(876) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(876))))  severity failure;
	assert RAM(877) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(877))))  severity failure;
	assert RAM(878) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(878))))  severity failure;
	assert RAM(879) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(879))))  severity failure;
	assert RAM(880) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(880))))  severity failure;
	assert RAM(881) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(881))))  severity failure;
	assert RAM(882) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(882))))  severity failure;
	assert RAM(883) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(883))))  severity failure;
	assert RAM(884) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(884))))  severity failure;
	assert RAM(885) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(885))))  severity failure;
	assert RAM(886) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(886))))  severity failure;
	assert RAM(887) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(887))))  severity failure;
	assert RAM(888) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(888))))  severity failure;
	assert RAM(889) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(889))))  severity failure;
	assert RAM(890) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(890))))  severity failure;
	assert RAM(891) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(891))))  severity failure;
	assert RAM(892) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(892))))  severity failure;
	assert RAM(893) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(893))))  severity failure;
	assert RAM(894) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(894))))  severity failure;
	assert RAM(895) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(895))))  severity failure;
	assert RAM(896) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(896))))  severity failure;
	assert RAM(897) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(897))))  severity failure;
	assert RAM(898) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(898))))  severity failure;
	assert RAM(899) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(899))))  severity failure;
	assert RAM(900) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(900))))  severity failure;
	assert RAM(901) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(901))))  severity failure;
	assert RAM(902) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(902))))  severity failure;
	assert RAM(903) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(903))))  severity failure;
	assert RAM(904) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(904))))  severity failure;
	assert RAM(905) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(905))))  severity failure;
	assert RAM(906) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(906))))  severity failure;
	assert RAM(907) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(907))))  severity failure;
	assert RAM(908) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(908))))  severity failure;
	assert RAM(909) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(909))))  severity failure;
	assert RAM(910) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(910))))  severity failure;
	assert RAM(911) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(911))))  severity failure;
	assert RAM(912) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(912))))  severity failure;
	assert RAM(913) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(913))))  severity failure;
	assert RAM(914) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(914))))  severity failure;
	assert RAM(915) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(915))))  severity failure;
	assert RAM(916) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(916))))  severity failure;
	assert RAM(917) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(917))))  severity failure;
	assert RAM(918) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(918))))  severity failure;
	assert RAM(919) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(919))))  severity failure;
	assert RAM(920) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(920))))  severity failure;
	assert RAM(921) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(921))))  severity failure;
	assert RAM(922) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(922))))  severity failure;
	assert RAM(923) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(923))))  severity failure;
	assert RAM(924) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(924))))  severity failure;
	assert RAM(925) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(925))))  severity failure;
	assert RAM(926) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(926))))  severity failure;
	assert RAM(927) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(927))))  severity failure;
	assert RAM(928) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(928))))  severity failure;
	assert RAM(929) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(929))))  severity failure;
	assert RAM(930) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(930))))  severity failure;
	assert RAM(931) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(931))))  severity failure;
	assert RAM(932) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(932))))  severity failure;
	assert RAM(933) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(933))))  severity failure;
	assert RAM(934) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(934))))  severity failure;
	assert RAM(935) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(935))))  severity failure;
	assert RAM(936) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(936))))  severity failure;
	assert RAM(937) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(937))))  severity failure;
	assert RAM(938) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(938))))  severity failure;
	assert RAM(939) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(939))))  severity failure;
	assert RAM(940) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(940))))  severity failure;
	assert RAM(941) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(941))))  severity failure;
	assert RAM(942) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(942))))  severity failure;
	assert RAM(943) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(943))))  severity failure;
	assert RAM(944) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(944))))  severity failure;
	assert RAM(945) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(945))))  severity failure;
	assert RAM(946) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(946))))  severity failure;
	assert RAM(947) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(947))))  severity failure;
	assert RAM(948) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(948))))  severity failure;
	assert RAM(949) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(949))))  severity failure;
	assert RAM(950) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(950))))  severity failure;
	assert RAM(951) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(951))))  severity failure;
	assert RAM(952) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(952))))  severity failure;
	assert RAM(953) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(953))))  severity failure;
	assert RAM(954) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(954))))  severity failure;
	assert RAM(955) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(955))))  severity failure;
	assert RAM(956) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(956))))  severity failure;
	assert RAM(957) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(957))))  severity failure;
	assert RAM(958) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(958))))  severity failure;
	assert RAM(959) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(959))))  severity failure;
	assert RAM(960) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(960))))  severity failure;
	assert RAM(961) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(961))))  severity failure;
	assert RAM(962) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(962))))  severity failure;
	assert RAM(963) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(963))))  severity failure;
	assert RAM(964) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(964))))  severity failure;
	assert RAM(965) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(965))))  severity failure;
	assert RAM(966) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(966))))  severity failure;
	assert RAM(967) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(967))))  severity failure;
	assert RAM(968) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(968))))  severity failure;
	assert RAM(969) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(969))))  severity failure;
	assert RAM(970) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(970))))  severity failure;
	assert RAM(971) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(971))))  severity failure;
	assert RAM(972) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(972))))  severity failure;
	assert RAM(973) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(973))))  severity failure;
	assert RAM(974) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(974))))  severity failure;
	assert RAM(975) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(975))))  severity failure;
	assert RAM(976) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(976))))  severity failure;
	assert RAM(977) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(977))))  severity failure;
	assert RAM(978) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(978))))  severity failure;
	assert RAM(979) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(979))))  severity failure;
	assert RAM(980) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(980))))  severity failure;
	assert RAM(981) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(981))))  severity failure;
	assert RAM(982) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(982))))  severity failure;
	assert RAM(983) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(983))))  severity failure;
	assert RAM(984) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(984))))  severity failure;
	assert RAM(985) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(985))))  severity failure;
	assert RAM(986) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(986))))  severity failure;
	assert RAM(987) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(987))))  severity failure;
	assert RAM(988) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(988))))  severity failure;
	assert RAM(989) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(989))))  severity failure;
	assert RAM(990) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(990))))  severity failure;
	assert RAM(991) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(991))))  severity failure;
	assert RAM(992) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(992))))  severity failure;
	assert RAM(993) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(993))))  severity failure;
	assert RAM(994) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(994))))  severity failure;
	assert RAM(995) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(995))))  severity failure;
	assert RAM(996) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(996))))  severity failure;
	assert RAM(997) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(997))))  severity failure;
	assert RAM(998) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(998))))  severity failure;
	assert RAM(999) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(999))))  severity failure;
	assert RAM(1000) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(1000))))  severity failure;
	assert RAM(1001) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(1001))))  severity failure;
	assert RAM(1002) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(1002))))  severity failure;
	assert RAM(1003) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(1003))))  severity failure;
	assert RAM(1004) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(1004))))  severity failure;
	assert RAM(1005) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(1005))))  severity failure;
	assert RAM(1006) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(1006))))  severity failure;
	assert RAM(1007) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(1007))))  severity failure;
	assert RAM(1008) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(1008))))  severity failure;
	assert RAM(1009) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(1009))))  severity failure;
	assert RAM(1010) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(1010))))  severity failure;
	assert RAM(1011) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(1011))))  severity failure;
	assert RAM(1012) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(1012))))  severity failure;
	assert RAM(1013) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(1013))))  severity failure;
	assert RAM(1014) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(1014))))  severity failure;
	assert RAM(1015) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(1015))))  severity failure;
	assert RAM(1016) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(1016))))  severity failure;
	assert RAM(1017) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(1017))))  severity failure;
	assert RAM(1018) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(1018))))  severity failure;
	assert RAM(1019) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(1019))))  severity failure;
	assert RAM(1020) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(1020))))  severity failure;
	assert RAM(1021) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(1021))))  severity failure;
	assert RAM(1022) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(1022))))  severity failure;
	assert RAM(1023) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(1023))))  severity failure;
	assert RAM(1024) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(1024))))  severity failure;
	assert RAM(1025) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(1025))))  severity failure;
	assert RAM(1026) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(1026))))  severity failure;
	assert RAM(1027) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(1027))))  severity failure;
	assert RAM(1028) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(1028))))  severity failure;
	assert RAM(1029) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(1029))))  severity failure;
	assert RAM(1030) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(1030))))  severity failure;
	assert RAM(1031) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(1031))))  severity failure;
	assert RAM(1032) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(1032))))  severity failure;
	assert RAM(1033) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(1033))))  severity failure;
	assert RAM(1034) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(1034))))  severity failure;
	assert RAM(1035) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(1035))))  severity failure;
	assert RAM(1036) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(1036))))  severity failure;
	assert RAM(1037) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(1037))))  severity failure;
	assert RAM(1038) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(1038))))  severity failure;
	assert RAM(1039) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(1039))))  severity failure;
	assert RAM(1040) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(1040))))  severity failure;
	assert RAM(1041) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(1041))))  severity failure;
	assert RAM(1042) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(1042))))  severity failure;
	assert RAM(1043) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(1043))))  severity failure;
	assert RAM(1044) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(1044))))  severity failure;
	assert RAM(1045) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(1045))))  severity failure;
	assert RAM(1046) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(1046))))  severity failure;
	assert RAM(1047) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(1047))))  severity failure;
	assert RAM(1048) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(1048))))  severity failure;
	assert RAM(1049) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(1049))))  severity failure;
	assert RAM(1050) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(1050))))  severity failure;
	assert RAM(1051) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(1051))))  severity failure;
	assert RAM(1052) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(1052))))  severity failure;
	assert RAM(1053) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(1053))))  severity failure;
	assert RAM(1054) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(1054))))  severity failure;
	assert RAM(1055) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(1055))))  severity failure;
	assert RAM(1056) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(1056))))  severity failure;
	assert RAM(1057) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(1057))))  severity failure;
	assert RAM(1058) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(1058))))  severity failure;
	assert RAM(1059) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(1059))))  severity failure;
	assert RAM(1060) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(1060))))  severity failure;
	assert RAM(1061) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(1061))))  severity failure;
	assert RAM(1062) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(1062))))  severity failure;
	assert RAM(1063) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(1063))))  severity failure;
	assert RAM(1064) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(1064))))  severity failure;
	assert RAM(1065) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(1065))))  severity failure;
	assert RAM(1066) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(1066))))  severity failure;
	assert RAM(1067) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(1067))))  severity failure;
	assert RAM(1068) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(1068))))  severity failure;
	assert RAM(1069) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(1069))))  severity failure;
	assert RAM(1070) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(1070))))  severity failure;
	assert RAM(1071) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(1071))))  severity failure;
	assert RAM(1072) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(1072))))  severity failure;
	assert RAM(1073) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(1073))))  severity failure;
	assert RAM(1074) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(1074))))  severity failure;
	assert RAM(1075) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(1075))))  severity failure;
	assert RAM(1076) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(1076))))  severity failure;
	assert RAM(1077) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(1077))))  severity failure;
	assert RAM(1078) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(1078))))  severity failure;
	assert RAM(1079) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(1079))))  severity failure;
	assert RAM(1080) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(1080))))  severity failure;
	assert RAM(1081) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(1081))))  severity failure;
	assert RAM(1082) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(1082))))  severity failure;
	assert RAM(1083) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(1083))))  severity failure;
	assert RAM(1084) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(1084))))  severity failure;
	assert RAM(1085) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(1085))))  severity failure;
	assert RAM(1086) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(1086))))  severity failure;
	assert RAM(1087) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(1087))))  severity failure;
	assert RAM(1088) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(1088))))  severity failure;
	assert RAM(1089) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(1089))))  severity failure;
	assert RAM(1090) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(1090))))  severity failure;
	assert RAM(1091) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(1091))))  severity failure;
	assert RAM(1092) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(1092))))  severity failure;
	assert RAM(1093) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(1093))))  severity failure;
	assert RAM(1094) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(1094))))  severity failure;
	assert RAM(1095) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(1095))))  severity failure;
	assert RAM(1096) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(1096))))  severity failure;
	assert RAM(1097) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(1097))))  severity failure;
	assert RAM(1098) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(1098))))  severity failure;
	assert RAM(1099) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(1099))))  severity failure;
	assert RAM(1100) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(1100))))  severity failure;
	assert RAM(1101) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(1101))))  severity failure;
	assert RAM(1102) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(1102))))  severity failure;
	assert RAM(1103) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(1103))))  severity failure;
	assert RAM(1104) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(1104))))  severity failure;
	assert RAM(1105) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(1105))))  severity failure;
	assert RAM(1106) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(1106))))  severity failure;
	assert RAM(1107) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(1107))))  severity failure;
	assert RAM(1108) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(1108))))  severity failure;
	assert RAM(1109) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(1109))))  severity failure;
	assert RAM(1110) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(1110))))  severity failure;
	assert RAM(1111) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(1111))))  severity failure;
	assert RAM(1112) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(1112))))  severity failure;
	assert RAM(1113) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(1113))))  severity failure;
	assert RAM(1114) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(1114))))  severity failure;
	assert RAM(1115) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(1115))))  severity failure;
	assert RAM(1116) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(1116))))  severity failure;
	assert RAM(1117) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(1117))))  severity failure;
	assert RAM(1118) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(1118))))  severity failure;
	assert RAM(1119) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(1119))))  severity failure;
	assert RAM(1120) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(1120))))  severity failure;
	assert RAM(1121) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(1121))))  severity failure;
	assert RAM(1122) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(1122))))  severity failure;
	assert RAM(1123) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(1123))))  severity failure;
	assert RAM(1124) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(1124))))  severity failure;
	assert RAM(1125) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(1125))))  severity failure;
	assert RAM(1126) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(1126))))  severity failure;
	assert RAM(1127) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(1127))))  severity failure;
	assert RAM(1128) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(1128))))  severity failure;
	assert RAM(1129) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(1129))))  severity failure;
	assert RAM(1130) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(1130))))  severity failure;
	assert RAM(1131) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(1131))))  severity failure;
	assert RAM(1132) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(1132))))  severity failure;
	assert RAM(1133) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(1133))))  severity failure;
	assert RAM(1134) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(1134))))  severity failure;
	assert RAM(1135) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(1135))))  severity failure;
	assert RAM(1136) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(1136))))  severity failure;
	assert RAM(1137) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(1137))))  severity failure;
	assert RAM(1138) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(1138))))  severity failure;
	assert RAM(1139) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(1139))))  severity failure;
	assert RAM(1140) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(1140))))  severity failure;
	assert RAM(1141) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(1141))))  severity failure;
	assert RAM(1142) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(1142))))  severity failure;
	assert RAM(1143) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(1143))))  severity failure;
	assert RAM(1144) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(1144))))  severity failure;
	assert RAM(1145) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(1145))))  severity failure;
	assert RAM(1146) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(1146))))  severity failure;
	assert RAM(1147) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(1147))))  severity failure;
	assert RAM(1148) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(1148))))  severity failure;
	assert RAM(1149) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(1149))))  severity failure;
	assert RAM(1150) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(1150))))  severity failure;
	assert RAM(1151) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(1151))))  severity failure;
	assert RAM(1152) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(1152))))  severity failure;
	assert RAM(1153) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(1153))))  severity failure;
	assert RAM(1154) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(1154))))  severity failure;
	assert RAM(1155) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(1155))))  severity failure;
	assert RAM(1156) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(1156))))  severity failure;
	assert RAM(1157) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(1157))))  severity failure;
	assert RAM(1158) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(1158))))  severity failure;
	assert RAM(1159) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(1159))))  severity failure;
	assert RAM(1160) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(1160))))  severity failure;
	assert RAM(1161) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(1161))))  severity failure;
	assert RAM(1162) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(1162))))  severity failure;
	assert RAM(1163) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(1163))))  severity failure;
	assert RAM(1164) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(1164))))  severity failure;
	assert RAM(1165) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(1165))))  severity failure;
	assert RAM(1166) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(1166))))  severity failure;
	assert RAM(1167) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(1167))))  severity failure;
	assert RAM(1168) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(1168))))  severity failure;
	assert RAM(1169) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(1169))))  severity failure;
	assert RAM(1170) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(1170))))  severity failure;
	assert RAM(1171) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(1171))))  severity failure;
	assert RAM(1172) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(1172))))  severity failure;
	assert RAM(1173) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(1173))))  severity failure;
	assert RAM(1174) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(1174))))  severity failure;
	assert RAM(1175) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(1175))))  severity failure;
	assert RAM(1176) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(1176))))  severity failure;
	assert RAM(1177) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(1177))))  severity failure;
	assert RAM(1178) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(1178))))  severity failure;
	assert RAM(1179) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(1179))))  severity failure;
	assert RAM(1180) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(1180))))  severity failure;
	assert RAM(1181) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(1181))))  severity failure;
	assert RAM(1182) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(1182))))  severity failure;
	assert RAM(1183) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(1183))))  severity failure;
	assert RAM(1184) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(1184))))  severity failure;
	assert RAM(1185) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(1185))))  severity failure;
	assert RAM(1186) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(1186))))  severity failure;
	assert RAM(1187) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(1187))))  severity failure;
	assert RAM(1188) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(1188))))  severity failure;
	assert RAM(1189) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(1189))))  severity failure;
	assert RAM(1190) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(1190))))  severity failure;
	assert RAM(1191) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(1191))))  severity failure;
	assert RAM(1192) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(1192))))  severity failure;
	assert RAM(1193) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(1193))))  severity failure;
	assert RAM(1194) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(1194))))  severity failure;
	assert RAM(1195) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(1195))))  severity failure;
	assert RAM(1196) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(1196))))  severity failure;
	assert RAM(1197) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(1197))))  severity failure;
	assert RAM(1198) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(1198))))  severity failure;
	assert RAM(1199) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(1199))))  severity failure;
	assert RAM(1200) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(1200))))  severity failure;
	assert RAM(1201) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(1201))))  severity failure;
	assert RAM(1202) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(1202))))  severity failure;
	assert RAM(1203) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(1203))))  severity failure;
	assert RAM(1204) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(1204))))  severity failure;
	assert RAM(1205) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(1205))))  severity failure;
	assert RAM(1206) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(1206))))  severity failure;
	assert RAM(1207) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(1207))))  severity failure;
	assert RAM(1208) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(1208))))  severity failure;
	assert RAM(1209) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(1209))))  severity failure;
	assert RAM(1210) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(1210))))  severity failure;
	assert RAM(1211) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(1211))))  severity failure;
	assert RAM(1212) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(1212))))  severity failure;
	assert RAM(1213) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(1213))))  severity failure;
	assert RAM(1214) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(1214))))  severity failure;
	assert RAM(1215) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(1215))))  severity failure;
	assert RAM(1216) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(1216))))  severity failure;
	assert RAM(1217) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(1217))))  severity failure;
	assert RAM(1218) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(1218))))  severity failure;
	assert RAM(1219) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(1219))))  severity failure;
	assert RAM(1220) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(1220))))  severity failure;
	assert RAM(1221) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(1221))))  severity failure;
	assert RAM(1222) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(1222))))  severity failure;
	assert RAM(1223) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(1223))))  severity failure;
	assert RAM(1224) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(1224))))  severity failure;
	assert RAM(1225) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(1225))))  severity failure;
	assert RAM(1226) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(1226))))  severity failure;
	assert RAM(1227) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(1227))))  severity failure;
	assert RAM(1228) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(1228))))  severity failure;
	assert RAM(1229) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(1229))))  severity failure;
	assert RAM(1230) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(1230))))  severity failure;
	assert RAM(1231) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(1231))))  severity failure;
	assert RAM(1232) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(1232))))  severity failure;
	assert RAM(1233) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(1233))))  severity failure;
	assert RAM(1234) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(1234))))  severity failure;
	assert RAM(1235) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(1235))))  severity failure;
	assert RAM(1236) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(1236))))  severity failure;
	assert RAM(1237) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(1237))))  severity failure;
	assert RAM(1238) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(1238))))  severity failure;
	assert RAM(1239) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(1239))))  severity failure;
	assert RAM(1240) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(1240))))  severity failure;
	assert RAM(1241) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(1241))))  severity failure;
	assert RAM(1242) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(1242))))  severity failure;
	assert RAM(1243) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(1243))))  severity failure;
	assert RAM(1244) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(1244))))  severity failure;
	assert RAM(1245) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(1245))))  severity failure;
	assert RAM(1246) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(1246))))  severity failure;
	assert RAM(1247) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(1247))))  severity failure;
	assert RAM(1248) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(1248))))  severity failure;
	assert RAM(1249) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(1249))))  severity failure;
	assert RAM(1250) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(1250))))  severity failure;
	assert RAM(1251) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(1251))))  severity failure;
	assert RAM(1252) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(1252))))  severity failure;
	assert RAM(1253) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(1253))))  severity failure;
	assert RAM(1254) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(1254))))  severity failure;
	assert RAM(1255) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(1255))))  severity failure;
	assert RAM(1256) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(1256))))  severity failure;
	assert RAM(1257) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(1257))))  severity failure;
	assert RAM(1258) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(1258))))  severity failure;
	assert RAM(1259) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(1259))))  severity failure;
	assert RAM(1260) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(1260))))  severity failure;
	assert RAM(1261) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(1261))))  severity failure;
	assert RAM(1262) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(1262))))  severity failure;
	assert RAM(1263) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(1263))))  severity failure;
	assert RAM(1264) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(1264))))  severity failure;
	assert RAM(1265) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(1265))))  severity failure;
	assert RAM(1266) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(1266))))  severity failure;
	assert RAM(1267) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(1267))))  severity failure;
	assert RAM(1268) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(1268))))  severity failure;
	assert RAM(1269) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(1269))))  severity failure;
	assert RAM(1270) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(1270))))  severity failure;
	assert RAM(1271) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(1271))))  severity failure;
	assert RAM(1272) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(1272))))  severity failure;
	assert RAM(1273) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(1273))))  severity failure;
	assert RAM(1274) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(1274))))  severity failure;
	assert RAM(1275) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(1275))))  severity failure;
	assert RAM(1276) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(1276))))  severity failure;
	assert RAM(1277) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(1277))))  severity failure;

    assert false report "Simulation Ended! TEST PASSATO" severity failure;
end process test;

end projecttb; 


